-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rzi0NqMp10Qg338h8/pXGxmwBGmZfGeLrtEHhyVhDfC0hninPYDdTSU7fMi1KP44uCCHyxP4lhaS
xRONbWm8uLJOQHz0e3KDGHo16wGGal/7SQIdOUkhynGJqX/xDre43xdOaXyOg2PCiUOWkSUt14s9
UleWh22bSBAX72FDCojudgqnP0YzsqJM2guyNAoq+xl73K7ZFzwGN2pqOosbYMSRCS79j0jesCP+
A1vG/0AGurM/C4DDQbwDSWfxTPwaLHegJmbt9I/0ppCfle211K5/a7XKAiU008qJR9afXOEGEI/V
S+QyZyDdTjB4H9i9TakYwo8xRDcrEHCiKEjLRw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9712)
`protect data_block
vOt2ApmDvAzPuddK6FhWNvliyqUDhr9fcap+T3h9vcYrFJHDXzIzK0xCgP8wcrIFeViID9Ti3GhO
PbFH2rcs8PKvKBu7CFPvcSouCrPceTSzc24fbgVFE18s75eP5PKzJkvi4dJeAjsNyTe0BV78kFbc
YBDzNnxeVUBDR8vLHJLAKWBK41ksZTCMqFpAB8o4nnskfQ9yFXSpFhtksJicQ3pDNOiXdVCsOvr9
svGAAOsDbG3vPMShFI/gvdGdb//TCwvs3gZICExPcEUPoVj87qf7TLWKFhMm1a13QtuTy+v9DHsk
fFVY/zfnpH1jJQwMaDLFGJ+9F0Hn41tkE/RglmhJuTfqhxigj4n39urr0P9B1aU+G9JKVlK6kjys
ugrMdvoHLlUGbMTwA1RtuJOORq7aOQyiH3lyyYI8mdlGFBXYhRJ5TSHgB3emYIIC7CmBria1iZ7+
eGSsJsGzGOHOWb61By7RE2z5koCRgD9wA9RT9KQ2EJOScLnljp0Ej2OmeH88/7NTIsu1eNEiWyWY
TKhLNttQfsVoAvXyuxBCjs3YUWdk7kVRWmjqJ34PBSoCCWWhrca62DmftfY5qkIwRzo6j++8M2L9
qv8f+CgyKD03QEMWJW34SIaSN1lnTFYyT9GlrJZF+07O1RiI0WmoFOA630FwbjSG6U8Bqy8Z9mAi
p8ZYa8ZRp/ja0Wnisu7TDcww0lJqlsSU1YHlVE8B4J24gOEoFacnoFT/T9RJxS7aDoslL5Ognymx
r/xNQovY/psyYFqLwQX9UjOmB6yTguByGcRzZyJjXTRAroE6rxXRB9dAhimrA67Y1YPUZHvXMz07
PlJbxWLCueMKHKxwXgkvwoniyZ6G+eR8mmozHpG6f9JC2s2zJi+8Z+OlR1t4vkycEb1YTTkHNYCX
dypmjfrRA0J9vrWovegmyMcHSIlyFFu/djmtFoEPZcxKSZzxZGEqHe+/NhD/dS023e0nqA2jp/lt
Z3a+Cytb1O+1mtwhJd+LgIypo81oY4HF0LdzQpa57ZcHUBCUCXqMPtCkMKpLs2yuy6jEgBSxvTcA
iprv6fpaHqveLxV2ANh/uyPFMEMANZzASf1XFxIg0t+rfvCMhxe2bBJgbp0TLUNrBWNFxJmA3pMz
uyln1nj5yYW5D74KiwfEWBL+rOlaDCmQwNBSWgvCgvFd95nFRvvTlMOlOb7Ger50UvGRwInMsvpn
NkRR2HoWekf3LXg1bm6kCktV0JFEhUorh13MjztAJsBaXadhnUbQroo2T1qjXXKktkamYfsOrMet
4cvwQBqZ7CLSKiktKaxzwQvME1YwJImTM+93mMkqeCdlgR9In5GfvTZ5PEyqlacgyAj+dOrkLwLC
agpQh006A8estWVARoud/Gz4MBWuoirv2IdtV+BnTKHGn3C8Finxh5zkEzIDIOXND5lU5++8wSLt
CtvICgae1Xg9qiKdFsS0Pv9xbPgYZ6ZD8Y5GdRnU06YVXBD1l9CX4SBjpHZzgkG+XD+HVRuUmRL1
nEh+mF7jI755heNKfKsJ1uIdD6vfk8ITTReDmpZ2iV+bq/PTKnbKQmIib9IQfu9fnN8vosOGhmMG
qhSVCZXl4egs8VYzhaYrDothT4kZf5YQxOkHMNbWnXdqHyHTXYY3MlrirdkBxLERMLPsuPQMZK/c
hrL9sKj3ylUx8aCEWEwUP8y4Ys4YU14AcTedeL2pfAe5phebYBwBQ0EonqTv1a+Ih3hxq2mlMrB2
9EP7CFc4EBJ8In460Wxfrkv4b6pSRjHO2QQqdv2PN+lAglgHcgOrgG+qh/Jwa3BobKEUA2d+sXAA
QzoeA0ZXDj9xO5FgJeJUynqjTA9pfNBHQHkpZtYQWVCIL7id8uenyNURTQZuuJSGK6hBEneCAUh4
XbkO4POGEQEH1NSYglmb+sDi/+AaeU0sdwDgUtDlMdQUrCXjBOJwjWxkaYzh8yuITifKyjKP0TXV
pfbdZ0RRs9N7UFzScr49Z5XCksJRBLr6WjfjuHm+GN/OPIqdEUhFDWbaLe3vIzyXbpSAFNqRRcYp
PqD0A1FU+lnLnZgAYujYKKI9AY+r9iWOnLAiGMHz7xijTaU8OLMkcozsRv63M1Q883MFGLGL/Vn6
ooudNWSt7ItBzZMYJj6H0rfNvDmaW6Bpjy7x9ikfn2btUPyDz0FmLC2Gfmmf4zYLTDDijdamMLF1
NBcWcHSQkYTAfZemvcmsKVxqUiO7hDCjuCze1iW9BRLHBEYwFwRJGdh6CQqKq/tFRo2RyBUy2VfY
JtlI4SXFqWrcS8+Qt+c0pToUEnSJMFSCx5OGXUgtT5XBSOI/Eb/6XXnEXBGOxUv/OFv58xXdUDaz
5pRgx+vDY6F7UVA/izvnWI3xttHP1HAdlFMI7BvKgsCSXcDmgAP4WDyHtae2xOqDMvXM3ZyzsR7k
jYw8va/AslmNL2F4yhN9PCxdjFe0Bf2fjmdYZRvzYdCAfegZFl0BnBA6pBVogqADSHcKZZQ1kEWS
wb+yIYBGfty6LjBRJY9846SwJjIUPOM3w5JsWaOV3Eq+yUNF3kes0U3Kgy03FkT9t2l9xpXPYFvX
Psh2XDccTdJVXpVDgnrXGf1Dvq+Jsnx+mIN05b4WUu9SwdK6OhSZuuzCA9WgqbVAaJ23osfnc1YR
D2Qssfc+s8rovks20ZNtID/wQty7JoHbLeZMXMczG0S+KK741dAx83qsIUTuymSyXaITzwpUL+Mu
Njfh8ZGEhCQ8AwtiM4jW/6L3baoVgwxxTbDFehLwx4nfr51NFwcLIXkoI4CTy+aIqHYSZc3mVYNe
jza8RaRwR0fBZZ0hFEPsS9Vo2i/YTNjIvdVWADtajRrDg07HIHhTlyf15cAysAe0xkidYoIDUWEz
RWZkI/4YPn5sf1kg+EQbZe3GJFFzf7SN+qjd6DWhXCu0VKHIXvzwPuKPaHzZLd1Cw0/aE/ahZkQH
ZyhWHyApUa23Wdb+D1mq7BniyflomwDcU2TE+IIEPGoJVhgvELQWwvcqsxDtBWvwTsANkWUf/UCP
iZlgeewZNMklUwaVKrNc33NL66XDqpXTAakAdtC3DcxdEqdpMQwt2gOKDqPwEsA6NiJd7gkmBEaH
v2ZQkWIjuz3niHwIu3tr6YKD5CB4DUVXNzFQb2GavVcWD5pVNJpq7f92RdO3dfzXb0+hkrm81fql
jmxz1WOsROMl1Kfwill0OHbPlEdTpRdo1PLczqWk0I0b/VNp97ePuYfLAyb6QGHP+29ZQP4dIdOq
Ci/yziBzEUViCe7vQ1b9QGrs/VLLG6JYeSaBG4AZWp6yEXG0zQDXvIDZ+rduBukUwUDVzZBeV83+
KDtqzTW9EOV6ddbm8vMtcPyk9AHR56VFJ7rvczStUcM12SLYOotDnJXu9R78zK82b0KB1yXslm+J
t1xu9A746IHwuWY5r0SxGRUvb7aIv1oXALXEURlJAW0f7CHn6AKfgdjI6OgGUR4js2q1hcXgNgIf
spThXzTsbbYDBCrGV/V3qJe1vXhC+YcFvHi+oamL+ZJFL/0Be9LGmcG+ob5xv4mZUrjGAcJBlF7e
xW1toBXG1a9/DmiMbUdVH2kB9LdNm90lwY9saTEo+BnUdyQmaDHU/WdCWf4QGRrFGqWqIEwRy5O2
n20PByGaCd1Gg+jo7AHRzFKu/nJYBUKpYoCTrGITY5GGEdqC1oJV4Dt94gv1Aq24yg4grXcIye4j
niXxu9kZ5QZOGPoNnq6Qks3CZlfUlLg4FvXN1gFobSx+oySv9BfqX+rkk8zBxz/YIXUL9ngkZ0lp
kw2MAcqq6qKGhIJtWyHxAWdprHo6nRM5FJn7PyBNa86d3pN+cMXJxLNbeP121CxL1Of8Tqb+IL6z
EVnd5eWtchOp49uhaR7jjuLS1ELKIgFbqnIfBqeP/5oxSkgxlRWEr77rSBsiWCPfR0jGozqfocR1
/NWm29BNOvHuqBLMrUr7nNrv1VdxUI0uARGEqXzVslHFdBOGnWODE8/ZvD/e9LpiyNHH2gKthm8y
ipLWhrhUO8p4KvYh2qcibJamxx/d7uCOP33b+Fe+RUsB9NtwB72JZqpsujELRIheYNNAJS5O8bJZ
eF2a9LRkBhskU78JURmUMTb5ZBxMgejf6DJwgS0deYLNSeLGZm9cMaQRccfHfNNOHsLfkCe3C0tM
iTZQaTf8Sifg9w7or3s8Sk+bCEyQhx7l6lMVncaEhp+Gnpo/p5AkDFyPinD41yfdguiBRsrRxFg4
dpaCiib2BfPNzpydn+jviuxkiLsPMTdmq8XlBaZxboeYp5lYiQzmxeMoN4s3/ENfDo1BrLGVRoGb
mvIUF12zk+rM1LFy4p+X92owHVV9RrkWw6XLIl1Lq0Rjfmb2XdQDyRbabdcw4mtJmhW2dF+4SbuU
XAcDUIAc5uhNsUoGQZ18lwJGmmX7fny6Bp/EQov64mPBAaz4052/51zgTuRkf4GEy5L1ZfgGr8jg
5ldLJKcuzPrEB47BtZi7UeP0qAq3cDgW2OLUA2hk9x9y9DJ2xEe0uV5SA+7p+ytiK7yTthJ/2gXI
9ygAAsH+tvOcN5I5/SMiP7T3xpz02RstH5GpcilcHHZzCKm5hn04jmbDuAka8rvnmXImeFcpPNhm
E9tNWZX9F5D3LuoTlwRpifZbG0noKFFAQKnLwjL6OjRe0lpsjMKUeM076aNXNQldi/GLR8fiuUlN
xpotYO6f/r39ntUTKWxIiB9bf6WCc5Pm+Zob8SV7o3pElmJaju17e+GTFnu26v4j+WTRP20oq+Pp
8M3skAbGa+KJaUePUGz3efNtB7erlqYkkL9SoK88C5ftcPZvKy3SiWVRq0abtFrhxrmi13Vot1DS
tU0Xl+tz4PMqRYF5oXXQvrRZHN4p1CjSCDn3VwXgGr/7vQWDIj3ZdZZsCHUWkpohq5QfFaZ3jpp2
E7ZZo4Jvu8hY34dF/s5IKvmu9BLrxDkPrbUsoj5IUzYpJFlL2g4NmJoFUP4+fqqJoqlnxRgzXzlu
2f09yU/OqabvLOLYBPYT5jctCyqz/UP+9iv12tjX+9YlCiYGO0MhsHUVhfZjFpLyQ4EHmU93Vdn2
hywKK7QlytoprRd270Ql5cL1FMOPfl6LGKXFv/lVuvlw7fv8TiDduAv256wXzCxLrqerYPejY5ND
VI1GTXhcpd4Bava2WVZhX6/k6JbcGmqwljIwQ6QMHLwW8ZTWpTbmBglRyTpGDLHjXzkgTgAtF3f5
45dnjYLIBK+0JwQVn+M2H/pgJY9o1+jHWt3kEsIHGxjgcBRxicNZz/fgXaoRMWww8515odZnyyhb
WWXWQAlp8hRrTwGFMkxJuGrprJNczji6fK+U1S8mxWyk+p4DZ8Boq+7rFvkohuxj7Q0T+MxQiT3S
/jR0EoYz3aWhv5VuS0W/LRrlMhMLM2VclSBNBdf6bMcARGJ8KQhZlesdy1Nm/tk2gNanoERVIQNX
fMC+cqbHAqQ6hq7eQN7i1a7Db33YWlyIAdvYfqR51dH17w7aUirFd1P//0c0my2cIEBgYgVxBUza
dQbEHVkjFjmLkP0dkJQP516uw90/qKMvgZ49lMZpTt1v+iFgky3WquZv0CFsvEKKBHqr2Jc2cGp3
9g3ph3hacaIEsX2dVAtCZrAVianL76EZVlwA9yOjkuBFdZVQ8V9mxQWPj5m6EojQAoQGS1BdmQ2c
2IM5BMD7VzghSkChyI6gMfphyRaHZ9H32yS2bNhYza7aJZyoBD+8KaI63O+FVtBCz1vnbqUdtliE
ATss7UCQBh4cwk+v0YdYMfveiioxlFx44+fvs1IsjJUt9ABzb/gys0niM4RMSBwbOCQHk5wqyQCN
yvKhGOWvdle9DHr/nVQ4tX6CDG0ZTdk94FJ8jOZOwDrVgoylF7ed8IzDnB3HA5oV6OwstMU56coc
guvRfRY5W7Isa8aHVrrIIIGLtr0rcK5XQ+n4FQ4xwvSMEsqaOgRzrzkdmlok+T0XbBBLUaZO6QTa
UPWMcr53O4VXYsrMb+AruNElAs7LfCPYHBxYn4wlyVKpIDwgJpBsSNpdBTw89YL9CYiq/D8aeZNX
5vD67S1qrAhVA8M7hRPDOfxaOYo/e0V8Ykbzz0SAKNuUwhRMckY37Vs011NpeT4WNYA2kgkahy8Q
BEfIxN+IRFLIt2JEBtjZHMgEkeyAGaPVR5eoVz5S0kg952OOylaBXUbM6n8RsAxspSwt47cOco7i
ztk9lqw5ePDkrADzXiNZEdBaQvlGfSZIFmc1CgpRbOsykxaCLkZh/VRoV4qEjxCF7RV8TmWbVciV
GvxxhieepdQDJ9HjYfAZfzoOAs75JgApc8lYaisqCIaZF6G5HWBtTJ1YbXpMhUWzSI5gLG9AGl24
nWdgMT9j46CLxFNATHHFtSe8mc9j2wOIjP0sr81qO7ZVtqvmAfDgNmIZFby+/3Y/f15Eit9d+6AM
Szk8hIiM9tvcO7FR0XXLtoUQ5m44LNsDzUWPStfpoXSj6VCvAEd3PiyAISlVs6YqEoSrjAz68uzM
3oRwBiHZmNTHDk3Q1Ru/wAQ41+z+oI3sXcfVtyRHeiXYAmCwLsMTStUU3skObipqaJI3HAFaCKM3
Kw5fVoy3cQ5rbqGboD5KDz1e0pQfXFh2GH5Oxr2BKbN3uvdtJcIhljWz87rGfxj5KwBJ/bdkfJ2Y
tTiucPbqnEXYwrF8dpn/YuRl5pqGUL3qChL7cjFFU9XEiLLe9jyDJDr6bnyfrrRWGNYBoyet6KjO
zCvWIBY+9KoSwIBfvYorqZi7GQ1RBI2L/U/1gYoljs7zGqmuHWNEpjpetVEwtYsMn7SHTam7EuY2
oPXGPN8x6ZW7+DR1kS4I+C0zuS0UVWLOwGJGKbgP4FPG5bTfCptobUbGUM8SHXWUVBMH2xfRodjR
kFySFd77P5TZMfMoPL9ixWs0eLmFu7bs0zx+Lkbv1KQ8WxOouT/cv0RChdWgLID9DXtUAZv237C+
DZuc7bS3EclwuYaAWz7vUUXLQelNQNQsvURA8mBxdMiEcYiR0Dp9rhm6RBsiqQYSG0AtLQavRPPi
zZaAqDCQjKrXJ7/fXh73quJDi+fOhPeGQN7uZUOy6ibW+9AAmhkuAc3XNQaxXi0uUFzKiH1HCsU1
evob6mguPbff0xWeibTy1XpAmj1jNe9Ojmm0+ON6misvC2aj2DkQAVlRzSgVnwoItP4WxIrFvjyg
2jbTxZzoTyvNaXKwxmBkwQZPtz3M49v/aHdoPj5pktfuTNXaUGDIDDIQBtHpY9PWMjyXMpQ5MFfJ
c3hwi2JiXS4nTKKslRqewJUkYVw1CqFqNHooEv48YRvVExTrnU4YxTvUqcZpkyXcAdVaJRyMWnrK
2WcPhtnuPc20VqBTIT17k3U79MmJpW5vza8oEES6nBVItvqLpyT3mzPMIwZb8kdPtrMQ78bI7AsK
L3mzpC8q6mO7cu/qHPmb+fzm/jWZRDh35Nijbsy39WCx2FHaEyUjmytILSWmaCjtWcY4pUi5HRek
hyBhM5VChAiObdSfqMVHZaRMhn1s4OQJWfokMl6apYbGmBaAxjNi5JCMe1Xj8LDmS8a0Z32fiJEw
anojgNAFQNV5/mmo8l+zKukV5MtIY2K7pE1ssJJSGlEPraE9ItTSJpcd1AoKvvwDVHBioS+KG9JY
dG4aIhmBb08vyYVqSR3cR9fqSdqOyxFkyOhne+EBdg0rbY63G5R62guwR9EjiZp6qAYQ4ejcf68R
44jONBP54CiAqvfBXw24WuR1H1Ui92l/JhefFgGDY1747ekYO48z74SoNtLBUu8Jc7F3ycbJUP+/
RLWC6HlFEdCtEW0Enx3ILyxcLShvKfXq/VKC39NYIQPuhBVbyGozjyB7sooHh2EqpCSvmWLr5x6+
mpYVzFcSVbtfkisTy2NjaqvnBEKFDh9DCSB5fFZBZOXN1za6jT+unQMqkHeSnvYBqzqx8DdQOE/k
sgNKESHrm7EP648mG4BIMnZ7tOcr73DIn12W2cjG50sLW/VvRR6o9qIesp5FpygOmHQNZXeJO4bQ
xj4a1kYFsceRwD3OWcVTNSLABrWU4DJbtfRIU+rq052fv898PVewBImhyDy4VN/QiXyqUsJcHfA1
29JsuMfZtVMs4ltg6kOskKbU1kkbTQDGbe8cuXqn5oJ1S3yu4LMnxYdRPZ4bldltTMGtCGCRjmW5
O79xLQ4gzcKIk13AldDcLY7eSjHJA1J3cIhjDwNfCvf2pKy6gkdsMTbcsExUJ+l3a/n6cwG1MDgn
mPc7h0OR1j6hpcQ0AxDkQMSEcgwSyvF5TZJECRToKq8QZ+yhHKctyhcmqJytkh7NaU1hejoMUpK2
uGP5PPPPOVDCw1Rc5TPZMpDeLOWh4Ln2IoN7bBC6/gU9EArKPYJYH9K5e0Izoe02cDkz6tGflViG
yK/5rUji9SU/ZMgIhp0H0UsDVHZHLLLTDwiCDZc2BLOzS5+wcohufNn3rbFGT7uboCzORQFiyuJY
aniJl9JefYW+RV4qp5rRZOvsPi5KQ6/z8LScfuz8IbM0h2LsRzVLnQbuAb3sE9fAyYFVuVHSIUZg
apxMIB9VuINpLNsIPpyraxAcbssHeo7KU4qDyfrqUXHY8ml3tBlUCPxbmkHxiXwtfRFcU0YUXuLJ
RlPHaRcG/jrmPO6Q2rZAjWADUGUjuCMcouoE8mU02UnYoH/FA7EJf6Stx9iIfzf1dGtu76unUM8V
952luFNhI0o2lsPaBdaCs93zLlytMzgpRkAC6hIh5VKCx5F0lHEXlCTTenFNVVJVj+0YpEwMUg1e
2VMCJcd7cwtrqVhsRbVj/69xF4S4NhsQFXqgzuzqjnqOP120PXkRTASt2EUPtINghRpqHg2aKfaQ
sU4PdT8wo4dDAW560mVBVNZo6ywAGLE4UzHa0Uxcc/kyuV46+doZzf088An01oSQFRwKH3Ya9Pfk
6vyONHF3NgEwcNw0apoDjgCk9NBocoLkc28fXHyV6xIhAi1hG5ZwC72qbc5sZVV8j/0FhksWMl7G
bywEFkkvvDhpIPAf+QOpIfQYmMtHwGy9+9HfJjdOp2ipn6KSWu3fkX7BMkh1+PO9B+EHP/3jBMzF
dbO+AOWHcTS60eLkMUa8Zi4Wb4JBKDWUbiAmwS8bN1r92cbZHzmoFfBZHo4s9lnO6gUm4YH5kqj5
HqFfqQ7fJbzfK7g5uczFXySwWwd85YcnHzVcMKC+LAVxrdk+PpUTEDJ+qxrnTeGanrrh7mk72xu8
+vXGTrDIMLNe7OEIcHgbr7p5thw9V2XbJuNBYaQCBwcXxjHL/EQKqMcXmqFUmOeFRNVhDsA3IA+e
fZotDTbXji9n/rcOww/0ALp7/QQbESZld/38GzDQ3UhfpuXl3LHue76bCiTVFj0ngil+pHd1G8qx
XCwWNWr+gBSpXgrUqHs7BENopO550O/720CaqMwlqbJtH35Ot5RVG+0nemqkeYQm214WkBQgvXLl
VgZ+rihKK1f+pjQjUtHRmGIsbPAN2JX7Lnba2gisvNAnvITO952RCZFzvWvHX1pf24Juor90ZFbR
z8ZMmmG+xdW3cUp088guD83NA102Ot1iahI1f+RbZFLN1PXChHNsZDwpbL2lY5y8inLqQTYFoi7o
ubYtXdtV/V30spAPWk+cADsMBE1zovDvAcJLPwO3ydZZOA5Je1l+wNV5rXie1ogCpi6Wbdbxyduw
NaowR1afBHaybLsxA7dpTZdZSmZF72CHYmyVxZ+4tPRDvX9i4OKtqpLMbWuJVplLask5YlcSK2/H
HjH/9m5aRydGKZvzjbhysGTjib9Nv8Dm7PeyJauM3WSd5MGzEseBclK5Dp+uAHfl8FRbmkJ0rblM
MEFrh0nfIy+h4lcDzMMGqEpzdUdWzcT6YoVjWcBjXBxokPENBiHQTrAyoxv6ljvEWBdzbHqwrpdx
5AX/Sf27LaS8hUR8lk2illLBpKzbdFTWsEzPavfrA6cprdbvSv9HayCCNByxLUIKc24g8pWOoBZ6
/s0ZDSmRpNMCYALDWftfe6fSY0yjpuo8uutM/YoPtfln/oorFixeeJe2cZGC4jGQw0LTGE50h5Q/
34Lo9tqkLZNLV61m2c79O9WjPzENbJQwL180yZESE+3nqpjOihIMV/qV8lXQ8yGejg0SwfMYBl8a
Ui8Y0+A/SN+VhlbDyS2pm3WyppsKbHlgrU70WlHzkrHarnNqFs/UBnS6ifDxE9CPxATqEWIzq6/h
kahMHEcj5q1L3skcGmpk9rFaCdj+srY0gBDwOtVKp1YTeOzW9WCxmvWWsEIrS77f6/SbBSpe1ug5
v/fNxJ2zJYxguUs2FpplNI0RphFfc9LEwRRYix2IhDugHk9YykFr1cy9r8hIZerCfyDLq+qaYVoX
2dkCGWj8OzAppZDp/ZEKaoaUP4tJvKI3s6wWfCGznalAqI0GOQE1Si/zX1EQxK+xYYKKpFTtiulH
njiMexD4Dkti6hfDc55ubpQOWOA93YGhWfplryRJs9McyW4gzuT04eUYDqLElDuKK59EWNmAStcP
TKThurcnRxoUyFP5+io7DdeAZE8l5DYa2R/FW/KJa97EnQBafQ9OZuSmW7ZZ/ohZo6pFrDbk87Qj
56MwRVO1IQB35IgxShP7Erev7XKs2vzVCW4HuR0ZHlb5qF6fESehavfXiwtgwsDo2mlUrnOGVqgM
83ZEatZkqfMP/Cf6SW45+VKwJJ5RX9BNfc+F8L50E3NxyhEwkWSCol6YOEFDkBy3RcMBJvIMXel9
dv/ioyJGAGAJtVhoebLkgbYjZLs9lDyEcOj/7bLZ2Tduss2sy4LGVVghVaNoa1HC6mAnFfHWJ0ZT
r7Bwfn2npqSVfEvcPyrjNOz5ljENnfDoMS+Zf7WPqN18yKrncN/ehx21P68zuaJm3zY6zNWnwW43
4gZt/Me9tg8F2SXWEe/3tfMh3C1fi0Ywf59t4t+nVe0dWdDyATD7NqS+e/io5RqFt2X2ZuVgDw/C
JpV1NPkZoGqMCcL6m1r4KuDQ6qiTfR6s8TcOsEZ36cbQQKkNAR/phGAsWEEqU4cMmfHHjy8SipL/
bVXOlH3YbBGGYHJjDFOGTBEb9f8M+PdKZnfGYy0URzcF2JV1jUBD8lq6581Hd5VfZEC0Ve9rWlle
3Zq+GbFkvcSq90HgDS/0UwOjCdmZIOOc3Z4yIR4jzA7uw/bEPru+8Rw7hcAax1LZLJz0DN1nbP+5
NCRTnmyXt3X13fIqB7itw2PpgWjs856WDEx+EY0eE97jqgDW9COaEPXJzsIE6WO5B0n7W0v6kgcA
MbXosVOWuji8debSV0J6K+LtOJq/AmIqVVGvQeQQp0vzepi7OJHxiPoKhSxDKKLTy5Dd+yHfeL65
qbNFH62p9AlUPYdDedWi0gtQgZnYJA+zceqX44XUVfRV7JSxJ6D9hcDklUUXG+VBQqCZguoTAht2
UlParxLSVzDr2eA7w2rs4tzCSx/rfgikecBPMtkFb5LJnQ0jaDsnC9Yg42LvuewA8O8BWidzP5Dh
bv5c0Q211a2hHr5ebBpExJqfU5h688fCJdHzwDHZS4Z3cL477x+k/dldvxjg1pPHF8lSNlqQvBhF
cnQctR77skpfv2kCQ5+yOuU+ASBMg8sTotp4QSckKQ3uZPXc1zujveueies6eSAXAIbySJTusYSi
K/a/AGbYZIuMF8/cVld1Heh+EAXsjaVUZLb03uy3evIU+n/nWc1IaofKvFOimmVyT438xxP8UTQD
kweG5oKlpw0NEB634mhy+U1mDnP0kzepDziPVPGmGgiGgFFZhQPYOrEZLJgl7OjEfuYTmboOWPu4
ONJV0iMFzQirye7LqzG7TKovdNd9A2Ef5fiBjFJxnYSJOwXYb2op6hjvbqgt1ru0yYx/B6SJ/35m
DRBWU+hgDKskQHq9/SoAl5SZlE92/rdT9OOCnkHnvVmvgrakzhp/eTMzixQosjPTelTjuVlYqsrU
do/n4Oeajzmd7rvc3pdza7Kemhfs057irv1LnYf3aP2O3XQRhNRaLDBFl0zWNUI3KaGhryiILwYO
HAXvssHMppjftcl7TQfKCb9ae7aVHM2Hm/hvXfjc3tW85gJIkE2+5M9gK0J1CG33kP5dxgMQ5a5x
qbfULx1vfMRJmowr7Bj7J3TDKzMIcEv+gEMTP35hdRv7um8NHi0iOLiM2sIz8frJ3rg8O6UJ0GgZ
caJA3JEaMQjNlYke89oNn6WQWGGxYL0WgOjW0R989x2yCy0G4hFNboOAWpgjpODhhQqPcUmk+8Ko
MYcEGzmMS+t1VTzWLY7zuzZc0tJXGxbm7kUYztAWPRWQJRbiwcfAuo5FZ9kHIYnrz6OZ69/GMbz/
FjmaDVYGHdI+jEcV8uKraYShRuga3n6zvvOZm3lkOrU0vdJm4lzIs0AGEH6VAoLJ1ji5LMAiHIC7
t2uT50ldzDRSVmd1blb1wheuWbXDTnmZZfWhfGwVj0/ZcOkFJpUrurWIEvtVy+mNtNBvMkbxj/Kz
yLgUbg4yoW5Z9EjiknETcTsW15CDGJFlhV3+CDW7NHUNin7NgZzrSHZ4kI23DoDO/54522jIPJMT
GyR9ucl0TVshJEnZs7TkH1AYSvT88wHAb/LqwoRUCbCUODwXlqj+Pf1u/aywAAxqlzQDJVmTZnPM
Rfc5NI9g16PENe73acxMXdsxGkacGVmj723vPbC1k//K7wogsjZau5TrZ2m4Emse4id/WJMZz3p7
jp2SDNO8+Sy9NnS2U+k2lTEoj720TIqIu/41YI7r18O04HuXyrhIF5/tBw/UpxXPZASAXK2LjfWY
yJRygu5eEocLdte4dmxzMUxQRrkB9PeZQ9n/Xjx0M6ihND2itSAR6OIfRRUz0xZ2t1Sqi1fDGY7F
IygFYv+XrgmGb0o8k1ih9pqNUkl/lA==
`protect end_protected
