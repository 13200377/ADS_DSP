-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
oDZyTy/+7m5NvjDTL+WklzAT8tiX7wMA7Q3QpXUfDynxak/grPJYtDcsriu8z9YNx2myzb3UDibj
ONOHK5RgKIpUJdbTB9nKnRIITAhADlpaY0WFglf+AhrACRDpzqyMHVRGbp5+mA7t/pR9y0owv5QQ
csWtUDX1jp/ihT88L9MvlDuDAH5FikHuz4yBM/WOus/kou+L3p/iNH6DVEKieN2PyYNVijNmahY8
yON7bbsZ+UXk2+VuuefSnavWHPP5R2qvPwBh9Bn096gIEe2TtBeE1ICvbXCs2aECaLMuzwMfUWqV
BQl5q7nFC40ASN9HdO+fD/g/KumfVz66l/xuNw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23248)
`protect data_block
m2JYUTXa8yQYZZT46DkNUD+FxTQO9We2bFje6Xt4Ns26OhAy3Vibd0L1ew/VRHtpS2ccMWj5tXZR
eKYwiZWexC2B8Zf6RyLBJ4oFj93XMqkWqGAtIneLXWsdmUQ9DCqAzsKuft626M4GXhgGz3kFLGqZ
Z/AvGdJqDEqTFv6o365k5pwm8ZOsX+KzwgfCXJFdVxVX3EhkKN21qxINPWu7fET5GDVcIS80YZyG
LS08aUs0x0UsiguOZTdfS+hDMkVqALYxfF5/xHyl0g8eZbygmS9/lhS03NpAEpY/4KbgAeszcDbx
3qr/hbvHtXfvxLdOHT+vhTzcY2CiQLslZgvEGnZWqxNkznZfI6DqR+LiCLWmwWb1txbTIjWL9vS5
4MfZTp58ItODei7H85AxycfGvzS9zUw1gu4Nu6dV//MFng1ns5IsMKMhiFfCa2X774k9DLsTG/Qw
/ubReIzE2xWtVfYHbAP5BUapRNBG/2fa9lq2ED6WUrkOpnwfN8RVjZ9asqDx5tTcTxY5NXFHgUY0
Xpic5rZE6dxx59eC35/uLjCAxesQriv3MxyaXUqFpRKUwE2GL9dCqIp13/rqwy37hWhXXIPpHnCF
97y2A0BK1L9mA/pNRPl8ckMwLxOujlkpjm5Y3iZ/+hFUWePMlh4C/AkMLjBLFTy6224gSw8D+FT9
OrgiqMxv7LJ9NZKyDNAd4Q4o36oX6dwlKWWyJ3ao+GYPS4zYNqkOV9H0fGaZzSrjmuBPviS5zANX
X946ZTQ5W6hvVFiwq72Pj0TzGQBB6DkRxbMAg8QQhKfFD7PVlGUUiXd53k2YhHJffcJWtXzybQ4X
SXFp7eRmX2/wsU4ZB/R//N92CoGhCMbup4Ptc1aEoJ6l2IJ2Bt0J0uoJABRI8RW5Edd5TeXh88vb
eb0xBsCaUHUL5z4Xls7ItYVdHRmGs/jqu0LsuJON6j3eaJsYDKm7O0Re0jCHAQckQquZ7Efq8+uE
tYYgRCbhdXlTCapjrdkOAQD4WuhjQ02HIvl3C7DOCKct21KgoKhvxc+yKL0f7jH5D/bSin041EmQ
9Xo5WVCVYGRv+iJ/nLlxujo12FhU0ojyzQ8gsRwdOgoowwNu9pak+YCkSquyOLB0hY6AEtHXGxGH
BVJDUaE06kY+HsN9rzWLVlr52YtROJBAlkXBJelVhSexYr9ks+MCDP213ys/euc5r1huS6K6nQJQ
nAAqBkRi6qINvimwduz6qnROJXs1rugXQ+93lkGfVh8QQw6voJnneG+W2Oi9bRbSkb1NNpURcLGn
gt+wz5LtVFSrd6sYZvFOaKYTI5qiAlRVrPbZCmgGbLbskFXGJdlUtWJF5wFGBP8DVsulWfpO0MiR
bhlyugZIxkpYcgXNeI5LHHlo1ACYmF+YiFr0Elfw86swfAoedGNcbRbOsTU/gNWcLkliGICFa5kY
6wvdGD7bgj6jXuaShKlH3+T6dpxfLBl3uXv3rhuficUSXfsiJGZhg1hiwqC4DMWedHxiBLEKEpOl
D6rG0RupX9sdNBAeix2dCk1gXm4Q+kRAB8xk4e6OZ1Wrul2xK1VpVLbDRTcUf1+OHhV4O75L5RsV
UWi7N/G4bcLXBniAp7UYDQzGfx0TFAbtUUedHbkxtyoOf2/K7DQ/BX4ivHAEXQrGPmIrmaqoB6BK
cxBYqqG7IqmEfXVcd00Jfm5ZYUU//2LQlSUYbluDx5YI8Xrl8zawttshhQLklgOlReUJgTg8aSim
PPW8+0TPIT9a0WkIhnKqx16FhCMNM5OjSs8JX40yxxX3dLzhY9TSzKKn2k4y8XYs5bp8NECpGbUA
1euUTxNQzHAnjEMTLKmFQahV5b8lDQPINWkOygG2SUj0TM5OjUc3OxKe/3Tomk4fzqs2dgpEtHuU
6tbg8cwfPmAmVPLbVRJC6aoDNBHfTlBqk6FkhSmZCdTcSn6w6faTGSNHftyO1bull1HE1ab8xXAm
wYT9XA21rdGPgEbXVvqllZI+lz0sQyZSefPSy2mKQFRYu2zfR1bELqq4hNAqDeDyz4rCGwQltctC
8jSzdImdFwooXlf0hGL5d2S7B4sxhegUvzK0y770AYn3pU0DjWxE1fCt2ADpBu2DvLFfVDjqyPjw
tlzd84+xBVMLndVJUAeJvCuv2qONPJ7ktkMpYWay9nit0Q942AKK35Q463mTeZAaJz9znL/+gfi0
J6c7yHwS47o4IhcgPSqnK917C0wU1raXHc1MpeTTA7jsZWsKGG1nAs7UeYaK8AAJ71zRIDLzYr6P
3FssuHXFB9soc2m9aZG4L1Z45+ZaSWPcGKI80+wpH+V1ECv7LMTIkI/7ReyxHmZtdJ+1e6rEKUhe
WJtkU0BcM/uOPxXXzsYDyrfyF+m84H1COlUIUf3+AfNKErpXJsdkhqVU4xn5Z68B4QH9H4PP909w
rtoL1TJFE6FoBD884LcjN41T9b0KWtR+PSyZskZXucXtPPkseF9PWcOLZmizOXstqMvl+9sg0MfY
kEC4VmOMPbAFUU9dpKP10HRUlM6l27Y2k2CEokC44j17WewfNsmT0nrHWrztt7W/v9pvBM4okjQI
i9Kt8DffxiYmxSG8Lof3j+yJIEXADC54I38i8ZSd7UZ3znOs06Qcfkx0yY0NCsFzMZD7D9Op0cdr
MUzTI5cNEEZ6aYW5e5EdFc0YM5JcdOf4LWBdos3EUlfTbJalv6QKF61yeW/bXnamtbaxqjq/iB07
m9yEJEWu+JCi+smIhgRisuDYv6TqdMu9KfXmCgyn0bFOFrzSS/9mNMPxImEXD2Mkn1kEKBrGqTQX
Gx8GeJU4sqjOprXsCJqADLSu4/I+nibO8r/558SNjl8T35Cxiymrfm4b86zVheli970fACDEKSFU
r9t7dF/4wZX9od3kdsKfzBf5Gj7Y788dqWrynx7APzCgtpb3bw/J5msR2YbIPS5hLa/VS4O8QOBF
k/zik2Z7c5ymh6jcduN7R+1ybFyS1fPIWULDK0Pkz0AuHKincBOcShSQ/N3BQ6WSXjegYwecwQDQ
VeFwSCus06GbEHQqt4Lug1mp/Nzk6AKK6ZYdTMZ1vMTEM2UL65a9bd6sRCSj2Ya2vpTsQqTl2TKP
t7vNgDA2aqOjqR0ed6mrEh7CZ1voPIJY0NqtjZNCmsH2EQSWBpHrBwvt63Cy4XI2reqlLazUp3sX
AGmNnfMgUa/zaEVSJX59s6nGGwh1CCiAhpHmSO0Lg1m3okxLvUMdl+6SCPP0xOpRyeWoT8DuHeLI
0cYErloJCCUIbJZRBFoVJ/gEY0ZBKdwi3FOUjkeOWxeUguttl2w7XqN5ZixFP370iWYGgdbYVCOo
RI9A0JH+n9LkK4y2ouJtlnMnBxib9B0rJFnwyuvjA8mw7rqZldza4tNF4PKAzdCpS2Bt2WdA+Otb
FWJSPkd3iM6YEiqfGFlqY9Mb3vd10Cp5u5g2+V3uPa/50qb8pLdQBl2OrU6f8Nah9FG7tFnBPNJu
1tGoN46oaJBvX3V6a25BdLfBeZ55s79M2+dEatE8rku8XOElFvSH9kb2PRwB3ON9OhgqO58o09E3
4oml+yvnJQCrJpH2Dbz16LDVhE9JNtzfUGiBNkHfK5cSkm84KrQGXW2sAxWZ+qFQECS/n6Tl8kcO
K0O4abGAJh2612xd6VSrE8vCHTJohDnZmdYUZWazq9tEtmd4b28G/J5FSRuYIkNnt43PWo/YieKr
4TCkFjzDbnUpFtVpzSAcPeVgtzOho5pjasr5kDQCzG/NM4JJaCEGcwuNzVzT/XIbaqR8fd7WlOZA
tPy4MCJ8YzPBr1wwb4Seqj1GxbZo5PB0e7JyPYRWvq2WQYRzPbe40Jn1Jie1qsZkQeEI9EMklep8
wI1N3Y3qmdWFf9qaRgWyhFVvVgYsAuXDcgyDajj4bxBXICBFaRIUAxQGWWpMErm81GMhEv7ktmnJ
jsB5TxK45KdJGl4HmEfT3Y37+Q98j9VsdysWziugsXwZJdy5ih4BW/2Wst5y1JFN8sPs5rBWCGjQ
iGvWAvGDNTWtna84aLF100ejrNSVbx4pG97/iw8eey0sONFUav0o/XynCPsVBvp5tSqFfIjl5efU
b/yo3gtEwy4DEl9SMCkCre2UN/hRJ7U7eS/R7ztKt2dypbexpnbs44S6dYgiQItERJyFmEjB7Ir2
bPbWkex7s2urvLA5PYB8kjJhAB2O5XbNc+Zw1J8ctiowurj1MsuBX/3Yod2i0J2ECWQUmnPkDfs7
7voDA6sBRaLV2HvbgQ8IgCPiUOu6TVHh16htBm61g+nSiBczBHog0sPG6eA9eAVkwKgweK6RuBPw
yBJ/zQMz+wwgsShmrq5N+muukvnPmmW6y+y3LYJEojtUKxAk64BjMWvIyM+wWWJwmbulcRRhIqBd
ApZdfu+NPFz7/C43NJRONAyP/P8CjXkrUNBH1VuKxAqDDFyA60heB/kPMAQ9015Fqqg4iUvIrhHS
Qe2jgKGl+gM64cQBHcbwT1Czz9hzf6PNa0QUQSQyi5YwLo0EvgGG1avJILoF+Vdc+N9HIpR5FTOB
OxyZr3aXraQzh4KVVV1jZ6wzYMoW2vvNFH2FQ9Jr82BsP7UiIQ274UpoA0zE4nmpncI3ToPk+IWn
CIvMra2Un4KxEBwJpkIwMwBflfiZz+uzVBEPphUDZwyHPVKKF6KbMY2+JnkcgHXE24AbvvSkrebU
t6pEZqK4XTRKGyGExy7GZcK+S2F7cOmY/KFAbymzK7Jsv6jTuVHgSgrLyb8tZ77xkJ4SStzu5pVJ
3mTnfLowxHHvJA5HXQDYLyKl6lB1yZiC/5OLBxOfLx7LzvOOGIGEveUH0E9gYcPCAhPoQXoI7fGf
Z1b2h/2SgNDCBnfMmiBLZ8zgLJGIt10m2LP4SER95TmKRNLQT4XL/Z/FOgXS6xzazY1lpYhiP4lA
4d7w5F+7rotIbHbwYBV0W2+MpDx1q/V15aX9gKqGkQrX+uQ7r/HByomzfcXqIuXIYDNdp4DMkoG/
zvDsC2tqOJoaEHo5HKtzDTabIVRvbPyFG8ctXw6iCxC6PxAgffgsmbwbP4z4RlNr5yAc7y/rPOvy
bkzm0aQIN8E4NDa6jCPAqV7ZqFIT83jgiO41bk2F9IXqu3YW0X5tI6z0COnIjRAvSy8y9UX7WsvV
w7qVJckz5EyNq02+Diusdq5Mnv/67dncYSZClFfDHrm5POmQjChu8epb8ND16kbGu278pbCNWd9P
7Kx5d9WUjPd4KvwjhUNkEGcahdT6chxtbB/iAgLHbnYzpES4h/8VfBV75HUZSfeCViLM1wkUIt3p
/1+Q1rekRXj5BuQTlz12IS2gImoBp7YzZZkVoL5pXkBX+he9u/qM8ytr/NA74HwqJCOXY/dP+YEO
clf21ASM/GLI6ju4gnoJveX5WPyh7IEZUF4P6hgfN+QVpeS+YUoPEInkknsKCP87ePevXQ4P5AIT
REhN0zFsB9P1Y/iYMyOsgNePiV0Dg1E2DOiBEGq2a4YEvCHOdvU4ltxPO2ya9E4gLpONixT+C6+r
afE7U9AWqiGkVVJrhZ98pLXK+Ba8X26VPIT6VBhgh2InDhsQ6x12pyBtO8AMzQhb6em7f4QcgB7f
akaZtCZo2v01J2bvCbUaexa8Ul29OB27iiXcJUZfVTZzXVodQQRhbXWpZ1VTk9r8bkw7qQM3stNd
Sqeumzody/WFG+YsdG1ctNJl2p38c18h+o83jn4AswTE9zErCuePQQmAOCES9P0EOMDj7BArE8Ju
LMeBFFulnPfDL7SMfyefyKQPfVWaEsCLt3lZ3rDoh6iP5p6D6vLJF7vDPE0gBrvXkz1XIWJP7tWg
SIcNWkKzkQHSUQ6Ihe44/r/uIm5yezjuuihpcDI+S+J9eTu5i3QOoRmSAk+mzCItktaJNx/ghRlU
Os5aneYm/kKAN5I5FcITEHDLt1QYHGtonWdwfwniVLwCTp1ksi4D0urjCWQaseb9uAM3BJwx1XGQ
EQxvZr2K613LHQ9QVsyBHY2ZsxQkDTAxkLdTsIDpVSYrTsGHyfUbSzoLq9DxRPmRSG7xpf/NlCYL
qekIUJUKwqQ/cRRFYRuU1R9Q2a5aZr1bilJplwZaNw239iZkJJR9ucfyKky+S/jIE7fsEXotGXhs
ZQxYsgkTkwrMOiuY9moQAecJTRaoZ/adc0ikKdGC/PgAFXtHnR/GEZKROWZcn2kHBo3QsrfS9xfu
k5zTXpwyWgMZ0u6LL1e4SofZZbvBjVRNhWid/Mgcskkiwsk92kmofKt+Z04kMS2kZoM+s71toIa1
UgLP6U6LLBT+VP6S/OIK7wM2e0rL15remY1Uv0EQtg0k/eQLYQ1lZldy0x1ZEZRTdH1N884eJpqW
beFldmRnQx0UaVkCfHe708D03fOePOmuxk94zDIqDfwPuxOY2jvrdS5AqQUMjjN4QtgLRUk9Yu/3
QOj2cTpYEPaW3Sb1ssFyHLbNWscpY6FAmn72K+oaRQaqPi5ZDiDuwVo1Mk4IIm/NpZQEhR2wdpl9
EfHEoAJBHqpZ7vsIlNPJ2B1ef9bFrmKlkzMT/axxjZ1FOHCCh63A4ynnwDvWcQbLOa0tkWL02Kjq
mEwA/rWz7DMaPCLqYr0ndyQ3lCBxybBRLKcsGvM7gRxFQm/jJ2XXa9uIEejDZq/pldJJ9E0SM4vR
cNGbjBiqXEVXWw9JNX5mOTuOSXTfGj73O8gSA8MNb9KT3lXekWYDgBy+Eyz6TR8Vn+InJY9Hh2G/
N+m0W4+vjmJXW+OOUy7LfOfaeA1PxhBFPLUUzOXJy9L9yeXZmaCpRnTAvPCpYlVsffPu4zd/Qxci
C1+VmK8tx4kJcbJOBKmKoOkvIZsA8Wa8RVmCMutvcPZqMF9sgPasKBqY47AyQwWSLXGWXlIi/E/l
Z+fFBv4xnS8HRE3Cu6vFO/Y2gRIPzsXzskp37mnyV4ptYgka6SHvcT+XAl8u09PbmGzjzY5Lo0ZA
3+YbqLARTWWTueI3JgEwjIs3yYH9DFnjtA4VaNCPkfgLXMFlzLrmbWlg6q9468v1IgAw5gWg7fI9
Y7aR3cbBXzstYhUELNrz7vnd8gtV04oQgHBCSRirrtyO5Rf9vroon13RTDEO3Cpg/VYGTVv1V0ac
kKDcnH60V+OsNOcBF0rtuSjALMha4VUljVKXExv7fMTnm719QAJ8RPKWF1JuZ9lBTtrMPZ2zSKT1
ItxghekPYTV89O84Gyt/Ovv9xwTa8ZPRaXtVUM05CiE9F2Jv5wCwMwLsk/OgYqEd4BY5OS3HpkbB
nJG6Q710llFRveA/XQui1NrpEMjM7lH0gUeRQlOj4KLRE4EQj2wS7guGWXhhy9LbtzT5a1wLz1Ux
Vs+S3ma+FyZiZai8cmZBLkZKIezqicPH0OVBqCUx9Gi/Ucl9s62SokOjxea67aDVu9NGyeQXoDos
36OIQl15cr75QaK32hoM0OYY+BQ5wR6c9xyeC3E14Znz9zaVgFfrnkOEJ/ZdxzPARhGr++ujNSdw
U9CbjJvSbZbmYFOo9/WmO4XdDhw6L4ZOLEA9YTs2n2XBzqrZS/Q/B8gRjNbiR1Ct/LYqMQuV+uYG
lr/lOLrONMVePWCPDoDOsbznysishIuagjO13DNQTGTL3wQ0QQvY1h0so+0BXNlq8NspzIkY0l8K
mYlR8o7u8053FXuJIB+8RS9Lmhfcpse/CV1xx+dVgBlKjUtue8GshpyuIjh9XrUQMOuR7EO5PXXM
tGX+blE5ths1sYZIAb9apggWH4+BnBqo9AjLKh8jbXPhpehngjglLHWdS47ekRxHXikuYHqxE6kM
DdbHH8qgyR/nnCakd/Ccqqs0Hokrv1IbZ+gQV4aYOVm7uoqyyaGhIb5ARtIb40kkbuLseXAPMdKW
/lRNCanThJAXfxFwJl+5XsF4odYl3+bqXkSCI+ZuMP1Ha61thQAMmm/TKjJrAW7Ra1U/WIbT9zxz
vvkL1zyFbEQRb7XGiJDtwJTpUcCkDnuGCTsuOepkx9mnxC9E8aS441xIV77pnBIUYis7zjpL0gbF
906pJaeEjSSNSQLIP5lPmcfMGcr/pyc5YcC1veyEIhZ8B9ip+yfYoyhj0R7Ztzz2qVLwklyIr65T
z3Iiu9cVSEVPPSUg5blSwzM5OIqHz0fG9+pmHVPAEOTZCUdJe7PC5p04MLBQIygluDt6HYQFu9CL
xiBr91alL3H/dpjOHLFrLzbODJlj8QaLi22PGIf9b+JVoKBhjUFN1iWf3daIjVgact4eCrMJV9TM
SooCzrl3yIMiHfUUToTKur4HTVACOj98JAR7ziQldwqUBVvd4bwC6bHXDe8VqBsCtnJAHas0ECKx
K1VdUFSgZRN1DgBlsXaEXj07M2XA/HoWjDp82seUP5kr3l59lve3g1Npab6BeP7kpbUrx5zZlBX0
fsxBPf8esI6eHAp8zgaKjR05HHRp6w3UcxyBEmpPOaz2E+cBeCstAxSD1YLgC13mvlss4ASh0gug
2gxjS9ThaLlVlFy6fGdGBbv6Zt0+LXwLVqktt0cEM5Hn5/tnIe53koAhETW2q2fQkzhwEQrbjflp
54PakeHt4MUAw5gdoHT+9Im1pgRXDx8WNegTxA4C5xnjMjYdXAIV+vYS3ZXC2hNmKngzYAJWH0ZW
rYwc4T54DqYMf/aWoPITyntJ3zKcVKZf8NKz2uHnfkWhlNN0U7ih8eVZIhB3ld9mXe8ohj7O5EWt
QkBEsZ7jRQgtPWCADpnCSbyBo9F92S/Mp3Jc+Ys+EFQqP0qIOSa4LMAripIZjw/ie1e21HE0zjCZ
h46dDjw1VMLBu4vnjz0+UTUaJwliJ1ccfL0HdLetkQG9jseWL8NpZxyom5Wt5yjV5OaN56XQ7Ygm
UvZ9JJXSZ6G+LHa7OPm1AY/UeaIzwcwYLLkyhScFUcjbTYAlu7wdeFYv3ndjR6kEcDgIBdfvpKIf
ClWdpoEEsTdawb8tM8/vKb/ut4Olaji0ecOTL5g3bN8wuGJ7yGN1TOBlNM22bDXmFKcQHTQoujLd
hWPwUX3TkhyvfFzJUNZ88TCUK9kBNzpLOV3WkkATBdKzBNOtoPA4b1Uj4tKgC+YD6KoaAvdVFD2J
Lhd/DaBhuDk5eVIwy3mMxmGwEYjX8SRd0YompQ6RMQ3LompFC5CXFIyxcp0BHhrg6xM7QcTa0LpB
KbctJ6I9icNLLY1XxyR6QH8cZTXu9gOPL8EYSXY7uqzPam3HslwVKCagPMsimI+kmZF/s9zFD9dj
F/s8EHda/RSGRM4T06Ox1sC7Rx3qTUrEFtPT0f7MiH2JXA3ezdeB0UrahrKEmwTZwS3jBc5ut7Qg
6YaiqyTElAnlHe6YbGEAIcNc5wcLaagtJoB7QkPh6sqPajr1CAsz0FM6Yui0uPmsGyUsU8PRAe59
jYsMEFF7o84ccOrJ2CE1YOx9zlPf1LZGxF0rT3tn1XBYCWbZCm2GT79QDyrPm0hDBZOaBJz4X7pu
jk4rM2Z9wdCnh5ftj5rS3QET+xq3Sbzc1CiaUT7JrHavppR1rDfhPck9itZ6Fv+mXNu4Guvs+amy
wGGu0o2a4LRlW+F6vLXkLaS6ll6RmB31MFGgAHSyeI8NysRloun9CC2mFS3rZpQHSvjZbNWToFEz
AUnIauEwYcqqfxqeBBkmJ+HRvtDWi5VBH4Cwu7xt03nuN/3TLUFON4he2Kx50gZdY0q5rtGslbQo
gp+P4u2nvd4pgU6q3eSJYPoMkKjE+sGq1pTBj8b3pCW7nA1KgCNSXbCc860tncxH077HvO1mvT+F
yT6edcwppzlwtXFKtn+awuhErfkaL/3WDGCY0LPpUtQEIflqo2BJCQyW6YpAqDlGsgOXea16MlyK
hYUdrmvM7cG/y5qHIpSg4Fmio/v08xMWFDtnfVfVXUBTlSsHAQlhgdxhby9FzowaGvCOgVSsrBME
01CFdHI6ny5Szsg5uHrJcc8A+5EhbJFAGgRCpJRph0KazoxftzxGya3b2A6xJZs9WdQun/JZ3Scx
mRLVR+QSLLtCbar6Y3vwc0LZbmRijLX0DeXdmAf7UzGVyVSDdo0foVp1C07WX8XgMWCQdQ7PNb1D
CUepCt25BquVhnB3CNe5KFIUSj6Wa9Ld01oo2invBNEvDQQGM8hK3SbRVt0UClfkXUpaXsRagnlM
OwQyKbav+KfRbGDhd/hfXGEMdcNs6yVWPzlQmz8gjD+PPHYsk/6X6xsOMNpBVT6vfTR45gDAbOuU
VvTVn90mmbGpZ41zreBa+MOoUOGFixMjSL7671j2hzFt6HFOJScSfQU+hwSPAyKxP9iQQrsjPx3/
h4/KAIL/XI98S24tkVxETIpwhJZURWTqPjryRMxvb9HDZxCL+sm8X1Y9Iksjq6aHem0az8wDeC+S
yRQOXcrpW78Z6j8fizGCkJcl4e+xnzIoO6LrBbcf5Of2wr4fP6Ynp6BYUL6heGTzLnieMyDaRdXG
yHx9P/9ihli+Nqx5pqwbbGQl5dzE0T0o0IVhnF3luuSnOuzE8SCginusSAvJtfg6ZeB/VHCKDCcj
Y6L/Vsxbvn35HIYXRHXXmdmDbyd5Uwn93xdXoQ+bO8C6i3tjpVk7yMqgyrAB8Zde+ArBofaPSjdM
Kx8f4v9I1y/6xlCZxI/xAgmLguadNCggsEbn/dE7ZfSTBciyEn66MNNztl80+mc2IUzTwtU32C+z
9Ftc4a0HdeEFTRUR8M5CZwo1oOzVGTIUlhGTds+uUeQxZATAq9XhZNUt3b1IIOmXIiThefGQ0aVJ
JgjUgWNN7U+/K4bvsZ6U/Kddu2LM0amwmfdaU9ilcHLocXZowuXWUCgRPo1C1oJbdTHK3MlpFYs7
8uMbpVpA+PfgKSGmjVB9zM6A4WnCg5MsH4aBEwhyHITU3RiLdNZP0BC7iFWZVOUZBg0F7Iw+Spxi
tuhUiKB/kWZhIw1jwgOf0CDCMqQGRUxgHLtiyPmc3CKNSgJr5MwX5f7EkqFiwM+KBAZcIVHAe4rY
TxIxRPpwUJeCBTZsOod5cncK9T8VR917fnFQ4Yugq929vWNITOZvoV+Uz2nTIRET5w1wzmvevWBg
jSHvSfadUc8ks1DhuKNgIcuCPQ1BolPyUF4MPWDtXmHd4lhP1ckVNZ6MUelE+GlQwzUz26e1AcTu
vksmXuxj8cCC0XE6smbOYpfOk3KcgwSbsC8aXDmA9OIQ0vkgzeMl5eVjG4cXSpozctROmR3SprIM
53PhE+zrOTC+xdlSQomz+DNVSXySKHcBwL2N0uULZ2fMUikXIuDRp00LHQOSSyHfxAvFfK2O2+TR
w8jICyrP9kpC1yOSS6oTLpI0LEU/sEd5nn7p9CARI1DrACoIX99lvU9jZcwaKfh+TIBtypN+Fc9v
nqld3fDKbe7w2uJ9j3WMFnPGfKmf01/3tEF1I42BYvPEtBuZtjnUoFcd2TkPoln33EPiZzH3UweE
ufyco9q3EkZLT1nu53Y8JFJjjXBuyGW3cKl3WIa01DRejquqhOsVQ+ewrrTe40+yjsyRm8kP5zcN
cB63H3iPJWIeKGRqZy2UHATTZOqRTU/nrTXpAXTJi3zFnm3LKtnMj8wH2deN4aZqD9CFeO2JTrtg
MPJrKEV2hsjc3i43gT/KDmiwJrNLiiILmc5WElWuu01me4kU6hkxPbjd8GxissEewvFB+BpmZ5em
rS6Ohn2jp0AvViqZRQyy/49Aa4Y5lRQUoPU6c9+2TnJsDyvmWwlrgx23sA/yOp6CcLCa3aM7M4AW
KRQDORPORpx3dXIvVI7bz72NofoeQRvKRnfkZHwGVwZcH3Jqjmjl9SEKx56r9nNRvOZX/DZa/FAE
Ka3KK6lUDJvLMpehRgzwNKvHS7HWEXK6Mm+07fRUt0aCxP6V7uSzK51EybzpwgcU+wZP27o4oUPg
uMA4G43bb4yKwsut8sMkyexIrt268H0HVB6q9sPuoSggRtKu/DaWqyojlscSEw6hZVS6JIyrEyC1
UBGe0WN0pSNZa34ehYCtOtUKt0Ln+Z0KrzFgWtGJd5gDpI2zb7AMmhvQpJEjvkS/LdCSQBO1Valp
5j3HqqIxlMvGsCTMj4mOPahKSNJeeur67B8Z4q1PQBF1ar2SUR9yqTx9TwuHh24Rq7ufxnreseWI
f0nOksYrsFjF2asYhqbqGcCQxh9JteGIzq1uWsMSxlfn+X+sgTyaWk7LvStsMDr5rLSKbOhysS29
vToRRijZN971p7C102RxIkPEFy0if9ugDMMPmpthVDCi6VZDVhKMfNc/2DDCZHwe2ygasziFsorx
E2ZR6XsKlSgfof032FcZAVJ0J4A7Qnilssp24gxNcfAWRmkGuj7+yM6sOX9EzKmsEispNo9GXe2z
Y58x3kueuzEqxtrmtWS5sf1Si3MCA+zS9I64AdGCqDbIIj0g2zcvZax+m0dy0DShOscGIHGkzfhA
4/+i8870DrgY4DA9pcXNi6fwcJZr+jgRaXlrISF5T+dvvQgsJAtntxj8hhH+wh/ZPVUg/zKjSwD+
J2KET+KVMf/8t1YPKld0NGyIjv9ynljlzU2aVdUA/PqE3L0SwubYQxn9dcp6jtv0EIhElAih/NUM
8IiqLlwuuGzK8MADESVP5UBopTg8/L+KXxJnpMOVXiGZmWG/exAMdAl+TY0r8BS2oTCfYgYmpgWH
P1UX9qcr04ogK5i8YaKm5Ba4lOFEOvjLZkqvtpH6VO+KwcSeFDgX5cNQshq+dToQy/5eFe3GgFLN
Vcr88a7TSKD16Kg3z02PLhtQc3brOW6qAsPpuottE6MxgbziwKicvF/nNTsKGdtuwFPQqvMRniOa
T1noboQvUU8uhhL0R/RcMJJlyo3au5WgNASaHQO3b17eEIGpvbVPbLIppQryNW+U6D3V2Vka5fpo
IwxtPNM/lp2z9Vgi6zgzXOtAkjsA8ttfBsVQruiijWokx4/rclixPaHxYlpY/d9p6AJFexhMTT5X
BY/Ownb7vgX6yKGY7lnGKwytyFlXbrGpb9QsfUHVeIqPpO6rkccrGlWN6ReJkLfP9dZ1OlgScw9L
oUB7vTnBaZomjebJkkVarPG5EOP0TYBtwTCSgcCZXHj0txlnSu3fxoxasCwpXn/4kXm3vI1Fhp50
yf1D28RAwukErRR/ycSf8MBR8hCx2BECHrlvHgYYI+e0gyo3YSuiqxbmud2vIkMesKbeWNWu4Kjb
lYMnQRqS643kLs5Db3LUST7PgcjctslKl0rV98ZfaZlCDnfh/J2oRqsG+lo3U2YYzqZbjgzkrd2J
csoxLhQws9pHkwjkk4Ii8FO75f1W9dKmq35c1hwE+A4YuQV04nGnPwGx5Rrq5mpbQZfOoM6rdxWt
9w0SR/sPWFqEdL/zNQSyFh0ZsKkTMR5VNik8qssI+qE4s5bODQSSh1HQTVE7k2TmoJp2ueLvBh2C
OufLkWLWwG/QmMFInfQDu6OfHINtmIc/OVjvNUCwaUmHRcJVCRr50hEkp9CXAEX6cIG6FkLrM9Hw
0y/EXYNXocVGOA8f4vMlREXXajUU7hImYP0ncpsdjujSE4OP5Q75fera5nrBp6gwdhCu6lcoAd6o
oyotRVUK2vx1LepBGbG4fp/oQNjgd0eFj3KF8ix7Ng7hGoBV0Jv4EGe1roPvTEJf4491S7qgeOaM
uWVyHji4mctO2W7c97O2hQBJz9heBVjEAwOraXBlr6X05k7yhVfYEd2BBnIB67YXPD2hT3NYuhxa
4IU4t3k18KGCJNJTaSzn8II5D4vUnKNdZdIV9GU2f6O7pF36QOAWXQMSApDiigMFi6OTFcRYyFwS
CTSrgTqI14aHW5NmxXLnOtcfYILSvEWFfm99RLETWrLdZ7L6cvRwRQ5IJnG+k4cYkvdWTIOnmdJx
WAN+kDEYwydL+/obXSQur/kgAKHoXO7nGenIzr6K2wK6/Mus8d1GuF0ojHVimOwzVGaoWn92woiB
+LgPhom9l8b4Cp7y96JvwP0QpfjEoZglAD1vHC3fBX2I1B++UdhfKV6Hd4jsanyggihpX1PH69bg
0pdVOit3bCKUEgtAGg5eOY5i4BeWDv1RoUJcZ5pBeyaiiK27bZOJoJV4GpxHWDuLv0KLO0+pjsjL
1coyjPcGvtfSROOVCP9ZG7EufapnIPfnbuvQn8YBWz5LIWdoToU3VxTPSmBMc/0g04QWx5FpgBBK
NpIyrwhLMneDpkZicRwRBP0x3A5vbpWdfqLuxhvcKrmhRm9U5W20k3n9qGW9Q5nCYwgdgmLMRUuk
p76i5AvN887ZVfRUpo8e+m78xyW+SQsBlz1RmUdGXEQBgloHRs5beXTgqhp8t3iRgtEy35490OFP
PgnQRHVseBxZHtzHtUOdlyMwcRHC6IxtleD8buVe8wa9kQGJzM/vCLfLwWqX5uf772+LcdW7lVXv
hMvlEeWOaOrWc32J6TQMqiGMg3ulry0IkRgUySWNZOVYPj0MegKXJVtICtuuolWEuNnftoe4JOXL
TNzwcx6Fg5pEsexUVw5241QmPy3tiIvhann/F2r1MXPjiyaQeK9+V0uiqKkv+ahQW7EwRf1l9VT3
4Pg/pAO1VgOx/rU7X7/UayzTRZHOFPxUzD2rDuQLJp0ZR/3ggCJyusYm4JzLoaOKC9ghvbRHRqWq
QPPSQG1IkJVEjvLvU+7vjv0YrNA3dp/TTFxAq9puu+1Ri+2oAeNfDSImhpcrpZ0WT8M7Qv+dXGbV
RGYxy98J8vtqQnz2YRlayL40RUeFr9BLjCK7BzovMeeUnAhrqwxOf08AM+KP2umyEqVOiNCJRKIH
sEqoHMVdjIGwa2frdJ1I4dPtgx8ZMnEn/RbvIatMowVFtBj4bvqxaqt4lY2ZuXlb/KcTx+koHh3R
wfAvVup+qGMigfEQsYGj4zwThMjEw2JAV+oBvinlvqRJtbENbtbFaqmrFhQBryvxUATLa80AkYms
1B3hBrxfLjGh8PZQ+hdElVpe92iAQgGR9ZTIo/Gbv1/fCdwhM79mqrL6YONciTWiFtHlIe/YDvMw
Z8CDGVWi85E22ReK3yZwZE72X+HNaCL0GfGZKeA4Zs00qNmK5w88Xi8DRIjsuKdqc4BBnW/UgdUV
A9MK8hLoMLEZ1I9L6dSG4o7+4rtH76P9S6h98EHBB6fkcl634s8alvNQsjUZLA/w085iYtVgB/uP
zl+iZiJiASsuTTwFTocPW4AkDAvYqxY5+hwXfbn1WkY+qLxq1d9cMaXgraj5BKtzwnCOkPS0sGV8
N7BEZgJ9n8hiBgsCQlzsW7QfYd4gq0bqdomXC+KWdbWpKXqw3HAAGD/l+tiZFwRHUasRrwb29ro/
y7gIjxW/fBia1ESRG8xKkpbCSUTUP36GJ9Bx1JFGUa9RSxgeCKn4+QcrS+ZkOTztBpIZ+/rD1xR6
aJFrNQMmI5UoDgI6RPfrfJcfmPyvH1UbkqjLE1oksVQlwDtVD9sgG57eLhRPYOn2hj4Tl0Wz7ryq
betHQDQXsRCWtGfyKghUOOGs4NbYiUNWvBgi0J7+iSApZxh/DfTuDtlHq606eO+tnvy9g87LizoP
IqF3qtRUAAg/aRQmUtkimPPqphjwEHYpHnruMV+DDovFX7trNeeWLMBZx9Iuk3XNWhv0r7t1ZsBF
z3xRBfPSzXYG/0nQdh3TyaDs2LVojwKzCf5LoFWzPRPPAf5Z6zrcDRNLHAA/UakSN21z5G6C4sAl
3+bOGYw4xriiqt69gr5VBgIvcgGv8sCklqwsImk1O6yidYR462I7aS2y2ZrKfgZtdvMMqycqrd3C
5eRC32BdvmPuqNyjrxRXbArYrMqwQBFoBWgKmk2ma2CW/+jGwKVukXXHKEmQP/HlopA4NpfCOg9O
FE/CGOtxXACSuhUvmkDofQSxBXMB2aSJgPFV68WOD+205EjadeIozN/anDPD32AA7NARbiRrS4gg
FMTkyTtNKqsam7clPYk1SAgTEztWDYyNUO5O2Wv7zcqkXnqMYluNUkxqaFEClbRPbOezxrBPPwA8
/bb5ihWNKxhUBQTycLMCOtFbi5CgA4igG9xYiAJgVn4IfrkBQCOp0yuwauyokXV87QznsQJ0B5ff
AdUayPZ7ehimZ3AyOCFBioBnD6dg1KckJsxf5D7KhRjTbGbFcHczEmvVx2ZjJqRh3QE8GO+MtuUL
7vOLKV8fFr9kvKpQqufJpR53y1ZhX/jSMcMb5FfAPixtXYQT74zmuWxDEJx/XwsdJ9HO7VJj7xDt
uszcAZlv45Kzg9spLkXKR9xSfvUCPBpR573mvqVALb8vNvQlNbct/d9rD0D6P0VFdma7Vbl2jcM/
UM7JKeMvUI+nKya0lcwtvfv1Xwi2ZLUH0KLIVjik57dv5SsI+fGiVfTaIjtffKUd3Z9/WiQVFtme
ZvgQO66BkBcUVoHViHJ3367vLcdNnvMrF+ik+I4KD2PPNCA21kpP1RbzwcsI2wGq/GJV6mVQerqE
BnHoYa+3eofP6dj3YDlHQXvtZ8P+CFqbZK/IMy6p8V9BvuLy40hyx0zoFfcLoTkYRs5dk5lUQLTq
63odryfZxz/Zc5ilcWoRrp/l6YQrwSLuIepJJCX995q0asJ6RyK2A/h6+NqBvZm6ofxKqLjz1yZR
mN9P82qJF/yB07tLbZknSE+y7YM0w9c3rGQAB1HFjLIEmZddRGDbAXVVI4jzxMnKGBLLW0zZiT7F
39cdCVHGTxpmBFD6lnkxhSZRnFtgSLZZSzL3M3wzqSqee6zHwHRXk0sm50n95gJO3+GSUPz8c6oA
zEwpG6aaA49S2zRqEbTuRWMvnSQy3rCG7HltKAFL60tji/3MtcAZCfNW3P+4KnT/4MOnREq12SjY
D2bISsQqS7tb192LoepmipICEPaxY3L482sF70ixPJYnnd0xcaveNGEmovilQW84RZiZbvAsrtrY
Sp+5sQSB4SzdCZ7TtgHSCNCJVxGFm8NvFcgrX6+AcDrrU/cfEMvuxOS/cUQJl/s5z2PhDkbmjQ+E
eGoNMVASqLUHfv7JVDyrJMSP6kaPcZyf1CeHlfBmawDYzzkeLf0aCQTCIYeMF1Gs+pkFTEtDJ9CM
717Wfaq8y2UsNJZ9mYc/GsUvAtwfj4oJ5jhFi5O7Hm2NmnyEeiqMNljft5VQUiXm0mgUHzmJTT3L
/VATeC1RAJYI/kMX4hqgIKX4v3eXrPeD1OxViqKhH68KlTNCcqJa3QFPMqwauc1GS4RC6nH90ERz
sB7FsgM81/Ys/QJyvgesjMcwN6lOyjJPu3oKjYVA9SsUa9XAMaEsOWIvgqa1hKtE/8WsVrGJo0me
gwekL85MXabNelF+UECEHhY8QYcvxkXsjunoAGlp++zBpJ8K38nadzZw7MLoZACl3grExHVqdT+l
/OqoehK4ZsNo+im7Mpyl3iNCgMeRi/+eIkshq8ViRUEawsZa9yGZtddbsmp/Y/K7uwKrxF7gTNR+
H4jLZGTXBfZLXXofZOuxC/Iy9YnfmvmJSQUl6j93hojN7W4rNx1LCQtKoVUcTW53cHRRXoPEYgrX
bg+CFvgFg99MfcEWJhNuzAA/0IkjciIX2YI0Wk/yvxYD0bk62rYqQq465hbsfDj4YghBFgminpnq
sLhPUSL7YE6yGak/WbytWUUIPIa89hvRWR1/9fwYxLa7VUZf2JSdUmW96BJLxvohSM0qa2jJ2q8O
uGdCJjG3Iea5xsIBhM0kyY7gmAbcIFGSl0xfJv31bxQyU/lKdBEuLe+Eo2n0K1lfp3+M2viuJ7LH
W9ZNWENLbvBx0cf6mF8NbiC/HPn0dFENm6SwQnUFA8S0c3qAL7v19r1AQC/7rj51peSThFOyUwkB
MoxS6sRGRFHZ948mCtZHERh8kb/lZRbbqeOfXityBrwG+O43v/eaAnvlOHwUiVZFjkPwgqRJZwwI
JWewWd8OXsDpMTccPtdMSHswddfI0krTEe5QB/SLI2d8lRseLozzWpfFyLpI2TpL4jrtgov+8Pn0
R6sgae/wJeUFENCihF73I0KRnTONtehkH+9pE0n7ydXwOu5Q5Pn3y3lajuuHDK6eqEYpDlGoDWUQ
qmFG2VYas8qbF19ARhl/iSAVeqgSvry/7XpkxTVitSgR3auo4DLK3I8V7p+SRUYp6wDDYHCtycNZ
XHXU3oqQ6KYwkIaSZBnDFhH3R+B6tFBzysz/2UwSMprK9BBBUnj66psYu7zZL2fLYPSNQbeO6ab7
18ssjcifUucz7vPf5WY6y07drjHfqOSfmEIRG5z7JbO+K4hg6yHFpuMtg5Q5uqlFZrQOBfu5Lxo9
hsBaBxLuoRrsk1LqRrDH8+Xs0efCriFGyojai/3BFn6lQxw7MAIz3p4AXisxeLO+TckU1tb0+XWF
iubhu3CeJ/rkhtGP9JBZL2rHVQwgMAzsOKHDnISmuuAMhAJCg9+cljqi4YZYZSeNTcsdVxTgN/VN
T706bfiGAWeXq4mCr71H7Vp09sDPPNtH8KRyzOyBDTEYDbibueusvhPsFqHVLvqDY8IleXXvaoZQ
+XD1lSLbQSZ5X6BOl01FQqxJFUm2ynyVOkdiFmk4ag6daYUmIPlCiwPQej4NexYE2hpII1X7y8g2
VnOdzlZ9LgHoRZYWcoYkOhdNgwMkRHjlC7ZPRoXIa7vNdYfmpKjdssm/24GDu5ZoU9ex5LIDMM4T
v37Enx7u6MZShzRWOKMxsSq2S3icQ64JaJllPy/afWL3sFQ2j4vcUMUIZsk4/g5FUkH1OhrOue3i
UpfEiJE6aSvsCBcABqgmiQtblXBByM1msTCEYIFK23idqm3+eTGuMfG1TO5pgfTf+2wWy8BwfH5z
7wr2Do5AC+ERcONWcxyibSo+zmg1/tR6GDUXGbX8aDxoDBPIR3CLO5Ytd9Fnq6ZzrqvNVvxEfnyA
Z6nmyQfFf7yMz7cVQXANsWdEfylWMRtoETQ3tkNbf8sxc+0wAyB+lbzP28ziaxgCGbXpiufz4XrR
CYiEzLyAjjbJtzRgYyyd/YoxLbs66gQQva2IqAgJ9skCvAVIRiP2jhmMD4z3Cc/mm6urv8Msd+35
HpOc5Rijudt7RRrg/JrJP5d9lzIQJT6u9jQxq5WtoMLpvdJUcHUAidiS5sUVT6Y2gvnnDLVbj22+
NLuXaO9WmCrPSAXcoyZhePtgbsT81lTdVEJ1aDSzUMNZDcfNGhMQ/AbQ7WvhrmzLYHBOotoLBs0D
k+FT8uWl4HZoEtzIMh86VGXHGYNYk4wdfoOfaXYCcUxAlqihAoQgUlmHKTVcsZSlPqzkTjo7FNIu
DDEyJ8Ea3EmXJICp9NXWV/yfeoMTE+WRXF7PheYeX70GI/Ay19gMlEN8Maqmg40tdqXN1oCXCKko
93sPvA8w3leLLvvkxpZxUZ6+R0e3ghFnrUx+V7F2xqgrf1oTHSDosHTKhAhzpqYH6NkjDTM0ycnu
ZOLvd6J1Zf9800AwbrVd6p6kaec51xJexbC4nSZAk+JKG0+nMZw43PeQfW/ZA59uXbK++p8ce8Ao
E9Qyk81vq/2cpaAO9o8RtyqQebYpBkJSw66A/BdJuZ4fVALP5Z9eo05aGASVb3leuYDxznvoPqhY
PbeACu3LomD6FnE5FHPTqF8/QCY9Tb4CR6b3LCXJizWbaoElRlg2scKt0pzCbIF1UFRSQknUScTN
p1JQ/gSy2rZ4np+vorDL+51DKq4iiY/t9MPSoZrKAW9Iflf/CKMsxcnRBdEvCnByyoP3Zo+iCX/F
WZq/JoWjrMimkO1spgUaHCedFFChJw1vDRwFcRE5xe0jShTEJ2OeSE2vakSac3tWsTRsjXog0oW4
Dd3rX3ybf5L3uLGsRTlRdGnr2gI61axmjd/ws+fwPcmNY+Sg6BdhAhgMBi6/0ZnKAcqiKG9y8+KW
X0d6vSdj2i6tPVM81FRYlffiSm+DUH+SS0fp9Srik6rm1XbfWtRum9b2MA5L/sL8EEMBmfg73ZPI
Rx9LVvWbBHm7GcAGXK5AnHrCzErYB7+2HdK/Nw9QYJM8azdzW3PKVL0r5u4/nK4sJ8o/duJyI2IV
v+IDXDfVlWu636GYpEgKmw8ZOuIrX4a/fCInpVzStIkZy/QW5cXSIuwX4Y6kEQIoSIjnMzRmb7RY
bV00nhcFodqg9wVPPu3UFyCfUBxZ1VJtg0YZDMRUTXWW7taYxvBRgALUcckblWorib4ITPcAwrcS
pSCQHhTu7yg07mF7OYQln3cj1f4thfxJWtXdVP70DvJM46VJFjmmOp59VrlsXBE9w2wlf7UO03P+
kZueJ6Rwumk5xwWIXv7P+MHzFq5Vri2tO17TWHMoMEBNZg6l1QcoHzkgSvZ54C1W3raTB0xjAjQo
lefglkGj8Sz4QTuu3yfiAXqZ+XcGZM8g1/JSCWAMWYXSljaXS05LWIy2eC2GcRuErcualgugDy2j
ZmShyC84I/c8V0Ow36HIvBFquBhpNVIecRK9wHAs6e5dObjCQ1q8ynu01mF8/hogyfFRU6rFqbHc
B3bz5yu608o3KzRZMYsXLlg+mCpn6hQHojI27grwrg7kinHJp8Wfc17m2Yffcguri0JH9a3uITs3
Uk7aI4HaPji/cyicRO8h/fsUnagW9atKNOh9PfZcIRxH4qzcNX6m208No3DRacPJUYAH+QUGewx6
MG9vznPszsBywgY/pZl/ojRIQ/RWmJdLQBkpouivKx8rAVzkhNg9LtzrcIgCBrHV64k4FanT1nDP
7a2TOrN5ph8QJoc+35NDPQWE18T0atifuTtG6L3mteKUR7AF7GIfUsOsQqgItS4lfY8GzzQFzp+j
w+b/QNixEu2GNMGgko3EfOg+4BOnC4gY0I4LHOZOYf3ouJg8cJ5Yn0I+ozny89vT5NJE6Gk3GhnG
hD4o+OHAP9TUImyNNd5+AOHlxnTfnpNMXYxDwEn4rlX+WtySZ9pQG/dTRz2JuakRsqmHtSII02Q6
IL4uaeJ5XjRQ23fOyGJd5MT28GPV2x8HsgxJwcKXUx+6s+KUhpd20WBVLe4/4ueej4/TnOtSzko0
SyBbUTCfk8RQp4kM9GlM6CTCAx6CVKiUhL0v7HBI4tFWTRhAmKVyZ63TSTUjg2487Z7cXmcqDKt+
CCBtWDQNKqmN3RdnFUfmih6CVP2vb0AUPbSwnxXQQuS4nR05lP4ETRncpI1Ovd/9aiTupdRy4CEE
vhEUf80oxKMlCQ7uyUJuAt1+oTEmCMOz2YEecms9dE2md/f0lutagKc07L6q6CmZ+jMP+9Cl8NNb
n8S9Y4qni+ykcboVv1CRIailpzCfA2gXOaIoQuDXIlsjl82+IOsV7Az7YjYjHej8oS6ldRet2dyF
+E8h79DzImcKwLSyP6Hk/fPOX/Bi3jgPEjxPjD8tLpFnTBeTKYoig9O0i0nMfB/bgJRg7EEXUHdt
z49pyq9o96yn7fcpLhUuyiPnilZ9ooXP8oedVNJi/JKE6dwzl4Z1puTIs0vV1do92qj1PduXosJF
Nxzoy/8CH3C7NW/V9GxK1HkkYnuFVz3x705PEVIgqH9y0wM4W/WAhZqe5F4L2hzQQu4X4OmscvBX
/toIFxORwMixAnmi50Jpl/X6ZBpoQ8YTjAMZh2rs6imd2DzuEjr67Vzh4bouMwK/yz2EBRdLqJn8
6FeIjtdIKbramAu4MhcVonxChJMCNxFfHHLyHvSOPvGL5nru2KXCycudE27FaA8yq2M5nfbhTs/j
trRFJ2w0MwAxJ7TJOaWtwoCVR1+7vH9j4Y58t9zgivvUttk8gNVgcLtxMYDnx1BFAQnZjZ1v96Wo
cerIq5uU8Zsn/8rnTCoXIcZZTNwFFw8ZV5xyMXXWMtiRn3SP874+/Wwa0s+NCkn5E2qkXA/VlSub
YPaIpx9afAfAASUZ1JBkNUaApl4kBJSezQwFDk6+UjtTWJ6iqoOt6in0g2U/tDKO3oOMctWEgSd5
CHHICK+9ERCG+uU1AbbHJ9LK6Mwu79utRDm+6jj1grKp4s1StZD/L+IxbAjBVi4g2/Y5j6/UbvOF
CpmZde1xmmGKfU8TVaMfZY4ZPu5KxJDPRvg8YpoyCfskUurFvxKJFAuF2hc5uVcQZ7kHiibcufIH
Jdu7NOJfyrqwOfGGha2nW743qDGiTFx5Ga9qX3rbzgpdrmdqwl/PhY267Tigkt3M+OfTBJJy315F
WqcUgGK27+5NdIolfgk82xExx8nZ9lkX/hGYrGpLj/eHWXJkBY1ibFnem8PMm/FqFZaNxQAp3q3V
bkk2khSrGEsnh3pCWWVNsHNuMMcp4BujkeGVuTcHLeaB+U5tyOuq8pru5Bsve5dPDtGkYmRSeQVJ
1UwYuwtfHp1B3xdw1NEOennPo10cQhyo7pcuf91GBKidD2Lu5cJb0LvLg5geJm6wQSaoKuJU6VFv
WCx1lXO2ZVAIS+k7C2eVe5c1xgig4XyupjCM1YpUaUhwhpFV/KqX+sMOskaUUF/zlRBbI7m8wH9w
sC6+2x5XpLd+Sz2iteQHE9/pBWcLSz2mp7I0llFszDioHzF1yWath7V521x9nvsG0+UNcU6E5fuK
Ad94TiEdBGj5c40RoZzgRluF2x1buRJHLc2CtJlM7W5RA+LfYvy/8XnO3iAPQkyOYiXP01M5zWMM
j6eXEMwSHqYer09XpFCumAmsGbnNrzyxpPM8hc4DJ2pwOz4rMEowpAnCRC8GORDiEGe2K0eJQ2DW
M8ZK5bRY4snVS4MEhV4jsSHG5ItPOvaY3InMhsPIsloMAny2xPlT9yP/RXJSh+HBkyA7h8TmBiQ5
SCJBSMx4MbBeDWYDMZSjdRlaIk0BH7bt2Eb8VQuBhwQ0UCEBQqDulMn/X3ng08iqS5HZsPSgnh+1
f6pmYeDFAayk1Fqwuzyg0Q5nQxkjyUgZmpedUWNNiIHv0CbT1l6xzeLWREScv3eMpoyB2x6N2PNJ
I5ijx0yddAMZL3sTXc+d72z2ECXOu2zVsFOO6IVHg+um/LhfmwXFWcZY0ApL5ZjiVJ1r7zc3cKGy
3/y/Q29dqVVL3+449Hx0rwyTw3vXtAX20JIHkTWbxDFvEwWtElKKKt23YiODCccciAWCXWb0ZhR4
3ADY1ONnIotq67HwYuXQkhEC3rCT7SsufYR40quRG2d/Bfp4fh0nomAg79awrtmLDRIgg09WBfXG
Mz4l9pvUYLAxBBtRGdNqYeX79o3ltEAxwXkoOC2HXNqCDX2BzsWzCbWdJvnTsmeKs9Ikqx95M3sj
FeNZ6oDr3L8iSgGrRs16QcWJpqFV8XOj4vskxIU9TKJoYrciAP/KXypXxAAnfAotCje8/r1h/32z
zhou1oO95HK2bkOd5RSKQq8BCuuQmEFNRhJ07GQhj92tDw+ExhVJG9cnn5maUcEkH9Mq8TqgGFAw
WXrqp47IoMdiPASnKvxDRVSP2EETeYtf2yBIK//wD5ZqT0QkcvMm5LrQUrG4f0gEgEUntS3Cy1g3
dL2RX40yYtNv+U3QCgU6itUekUyl+qQNuMXdqJyQCL23wR23j3LZAYHlYSgh7nkYbYUQm8uZim1C
QqHIOTaaTe2xJTSBYFE9sKFErGjJUfNk8wj5Fe1qLecFnmJqQqndLilpV67OER2Nvbe+UvHtL/gO
9k7DR7KTaDuT9A5gaLBmnxbPYb4fAvCvbxZCh9YbeZLqoO2/w3oxeyoo7LOU4ykm34Q3RpNLuhWQ
7zXbAZawpSRF8DfKvyfkoecHadIhuyAf5R2/UHr+iW/hUG1+MUVkk5mj3mP1JgjHc8Z0lmrKJWuZ
cbBc3XBkdzr6K9qTJSmpudeMPJl6jz3Lc8IepPu8WnnNdFrwdyE0sHOFyvfrBr0xtVxwCgXxdyMa
JlmJhCTC2LnhRUeoLIQ7IgqUKP+6EUdzGdk0SScCxTvW2rFkP02gYDVtXkFkGwxUDvq0n3WDs12w
WEzX5aEsKmvt3nvD4ycyz+fJ0IMqiF5Hn3BKHvr2GId22lyY5A1t76euhZJYx/STf4Xy7GZmhLWD
v9DlWXMqkxQ1qMZMiYBmrwEYghu8oGrV7Pk5I7nZkcje5/7pTC1f7fMS1I5KmW+CR33U2+8N9vSX
SEfJ3MEq9LTxaBZD0EAu2CX5aJ1DcxtynLsxqSlL+KR90OLE/ZLTGPteqEQtUOpVXzIkrf0E6LAM
7k3P1EI9pJlNIX3lTnxl7IvWwixHON+cr1q1TGZv7S7MK5SHkUY3QLLVQFRlzYQnlg1laVC68ijR
SppbQXymbNzBuSj2gHbrHAo6L24r1JR3kLSLkGU6ZNzwO9h0+zHovuG9cZmB8aoVmJkGgDiusWCO
TJ6V++mY+MHsCMY7w7M1g56wDjsU+nwQbndxxEGRfjuxjkfdHZNSt9BJwZLOjND8PnS4r4pdGPtG
dOaObvzPCzK+3TNYS+EokhRuBaPezh4rYBy3NazEqWk/FYzYHrceSwAen1slhcoSpHRpN76ZRgIS
LAl6rBryOkt9ufWH0i05lbp0DRnYnfav0hMiFON7U9cFfzhF7RsE8KqvL9ZRp/nhKHEGyMAhswAi
JcM6T8fIPYhQjt02Gz1EtgyWjrARM1lNO4MtCEljvdsoKR36axqhFTe+erSJs6i9dJ7SoJjvEEyW
baUH9G0JRQVxUwhGXmRP3MsXmrBBxb7cifnLreo6jDYkV6z0GVI7JajHVxNvLsTbNVonAqSXk0lp
Jnex/J14oPcZcbAYAEeyijlMBymBvWMo3k97xYcRtkGFqb3y9iHOMVVPEXhN9lVMgODJfq+2nQ0J
LlTZWoE5srMR+WEkHXXOn1RqjggVljVibkXg2tbj8nxNdEN3ULA46PFIePS5g+ucznaD1usHr4Ay
TAi7SNxxkIECr3sp+zpB7e0H0ErsNjMlh5R8pUrEEoRlUm6SSyw16G63kUu6LkvAYBDIGuDwKA9/
pgjq6V8G75Bm0cM7L+cfmUFrO54zic+WNPgbJ4PTZWvYTh2TxBniVb2N/3/pilzEE3g5/kqhs65y
+ZAy6w2UVA1Q4n1se/A4WywPfBinNiPxURN8sRlVnhdtACtlwGzrZIaGUyC8wNHmtS1bPsVnRSsv
iDgPqySNkdRCf+s9VQ5+2IgevTG84+TcrRjxD7VOzP56HZoG/AWNanFJ27jHnA7Mq2uMlgljkjLi
cBhl+lONnT0XgmSOqopEWf+Pq8GgTBMp4ta+4PM736GlPOUvWWZIydivo5YEc2qVEgS5hiXZ1PSX
0DfLHgUVeQ3pVOZD8PTacD/INFMWvgJQee2VlLKh5IbKKUSR4CglNRs4XYD3zOj8t8TIVrbHoPP4
LebeWwd6nYkKWjoFyoKPY/zuIBkZyQorWwqqp2+H3r8p87vJXvSS0Q0UfeZ3vvQsPO7iUFtLrp8p
wkwZUw8gdqzi6iJQzY05bOncT+8GxvsOvA2Z3EuspRDPF6zhQxJNyCoj5GU2rY8O7dbbshVkY/4k
CoWS4CJXUYQHU8erEkqOwJDmTID6XqCOXTzQHxzwOqz4pcjpVQxyCof9oNHWGqw60ALhbaTvnxgb
ybIQVZYCwKvzEF0/u+Co82MqL8IEAa0yi5GlYra5kyBTmvVuANfIvqDMWEkiqF5AJrFL6s6XwY2f
+bTtHRuBRt5CKWkTKoVZjw6ebczQzeI0a+8rynKZYBZIyuTCnYlAAJzhu4coXnPZjRRF35n9WYcK
1ErEjoPyiafUKxNRtRs1vdJZwHCCBuN/RQ2vJeXkyvGdv3NG8Skws3oEhGfdybEui7NW6rhd3u/l
WFWZ5I47tJD1lz3naEln2cNZpvNpD/P8qrWHkbMBxRqlXZ+EIvG3VeDIR4D0sM9RflWmlu2+Ow8k
MZhjCu49+VW64Ty50xnI4G42zX39VH5Mz0vWHb52t4BFBCHapH1EbYG+fGM2MW9RV6zw2mXbnwq8
PfUVe365jyNiHbzJOZnNQbGhDPD8/s43brQXfvR6nv29HoGVqRV+XHrCWbTg/ISD8CjhvLgsGuXm
44+q3a+of5LhtY88/HaPmk3Wsthx0+NR4UIehKVsvcwVof+wTu4aFYlKT3brS/y4DCnY04iZWIBG
J66uLR7kzrDWAg5BPK80PyCEzvQHfqFLbqb19/kYq2zaXQNt4RnNE2qI4M/po+NNUcIZA7t9jQtP
V8Qjlpb34fmrXdKMHbZQBQhZ8KssETaJXnSJH6iD7D4i3e7DC13t6rb9tYrx6OlKhtBzKUFNY/Pj
71AKYl+Umna4Y6BbF9tsQwqRijcze3hfifsBSEynvqe9nIwyWXGP1z/kKuB6FvOazXC0Djp14Ric
mho9WvyT+87TRt5C9oHwQeezcNSev9jShHAj6lfh2ObZlaf7VQ4uX9x05PbOQbTK8n8sYYg+MEmc
iUs57Clp/z2L+5MZYdopFZouGOIsgEeCo58gvNi8G3K8/cFC2Ja0BrBR9Ex3YOFGO2U18UaHOVqJ
lyGE0uJ8zHgkV6nTXq44hvCu+Q842S26HAdGAb8QyJxSpb2oonufKtP0bNbre1p6umSgy3GLx6Zn
i2AdPdiqsG+oGX9j+9usfg5J875JMjXZFJ6Aaiv6Y2L9fyMSx2tDREkA3cVSIj9ZuR5oPFLfi7wv
Oz+/sccdw4e4XpheAUJEBV0mCDJxKNrolEQgkRLjLGOc4drSzLgALAy+2r6tED1joIrL9CzaJO75
dpfAcU5OPshqktU/GNXV4YB10zerQ4U6elnqIWZDNTc7N1ZxsxI35EgzJL4wbO9EEA2HICfdaCrq
wvya6Bg48T995DrXVM6aEYa7EuzK0mxv4RH34hy3xrFOy8cbEfDUwdcWOus2+eIOyEONys/S8lMG
zRjnGoTtZf0ujyIhMv00QVRPMB5vdgggSa8EpmiZi3qyzw7b8JxzrnsktJCTBNGCNFzN5uKwnPlM
vVhYfWY32X23/BzI5zOqrVeAqlaiwA8GtTR90foGlWSOJBKJ3fImEHl20sblbZzCCtfYPVYuriEy
kWhsKgoaOuVAT0T0Ai9r2WIj3LGdhLoT2MMS4S9n098aqYBRwFkdmjeAXBh78P3z9Czkpwl6AOth
NI5GX5rDeNDK8622HYaMmFbmJvL5I5ZG8Npmi68bLHCHogMns5jCHC75vjwrSkj2I08B/+ao4jz0
VexHYbVUcmJnUfMxwElpisId8kkTBkcAMAz7bV8TBsM29Hbkvr3m1hilKy2Wxmx3UJNRLEc6JByY
cbLO7AlmXrLWHJcN2rYTp3Eh+Fy9N3ifJ6gaLIrxb3b+KFyRdQOHurErx3oDRlCQgvBxWQajlNYu
LY26zFmZsdIz+nQNZuPORFp+4sg5A0Pyr7OsS45Yyq5moZLzyhR3BUeyk42AWmPvbgvcwMR+yRFG
iIy8ISoMIl+r7jIcCxJirb1zzo5ZqPEGPpC1Ko5KKdMvW/lzkyszEBeAgVlEac3ex5JFrLpcrauJ
+iRgW6GglEqYfMCZ4dOvwJDoJqKKuDfn9pxqvWvdrrc3YcFmC04UHxHpiIdmmwQpFMvUVbTgHi5V
WmbCR2bYziL2z3QoaKLm584k+8fP6EVBg1x63Dfa+36bSPju0gKaY4wyed+wTkGNUDQVvt73zppd
vpa4MqNt3RyaAPpQ9ThhDdFWjpPfrPfj6Rpv7gnZnz8EexVx7tOGO8ZXxMiCQwlDGVhrwR60B+F6
eQtXh3J/gSMwwKEg535C2sLwYJ/Lre/AZvGjy9yKE2rO+NYj3dVZdwCxj6dseCs8HFJGXGbGI6Tb
HVZZF/EKF91BqYeHfx/kwu0PbNVhR1hNn92X6cLH7tidh1MvzESpywXZLYfJ7ICXV2EJekqWR7qG
q7TOePtxIaVoZCxt8lpQ6ZlxLQLfuH3xTpGMkpnhWv4l/5KfAXUsyQUviABk26GjQcCOZq02L/YW
ZDhgBGtglKlzJidk2BIbKzpo+Pz+vO1AlaCgQH2mVC76/lwEN/rwdoeOkvPOoiz+lnLGSszgy5Vu
bLieJC9J4N77vLKnavRYhOU/F4SecE1tMLADdLrw6I9DFkIiTQK0AHIR1UNUvS66Ec3eMUNqWXCx
+pg4++njnPNiZRU78KPqNLzZYKw0Iah9W/ULmuzF0tPJC6B/dsEF1hsc3W4nGh3YuiLY+8fsQUO2
9Ydr1v79vUliJWJVOrStFxIKJJPX/sjazj3t3/3eG9tmwOsr2VLKmQjZgfJKpnZG7y+OskOW9aR3
VVHfUIjBzA2vpgkJ/zxnnyjFBTkFbUI6YRhzjejc8arM7cGOZzGc2fe4v1+RioStJ53JKITW6O4Z
KahR+5C736ygZJ/AuTZdy2lpTaEIQ3OYx5dJ5LMxLH4z6cOkeD05xx2EmLV7w2nfETwDgugmL6Jp
v9hYLEEdemc15sOASjbN99Eeq06ALZlEF74zKSbC4sRtWdfH7vdMbySdKsPtfebrW9DbpRt9qJ7E
LHwiFtEXP9Iju+UOWXSQxT+woeyBdXfjZYVio1ui3N0lvqDu7wvFui0fjPi6kWVaduEpiALhPEYo
bfapgmRDoqbEufuPiFgzf+neWebHsTxagVo9sBBnvL5Io3UvS7MHRynKWe1MHczvZTobm1YIqpw/
6a6i2OZiIBqXGLyNtvzO+G/ZorImkQjSV/klp3hzszreeeewuifXnHw6R2YVwbgR/JZa+1KQwJf8
E7aE19YjQvg8b2N2EMefc9IIdBV1PKveuoV2IgGpeGqd6HRvNFFu6BK4YzlCTpP+/vC+/lguQ/gF
b5Q3tD7/aqcwSjeCjZsEnyyP/CIUCZqvJkZgBI6fbOuSMrfanfGFQU/0jxrLZda/6wnq2P11yvHZ
QCjI4GPRwgDdjbtUAhWJtBkzZw/kxTdJSkcEoEFGgtHaTSztCuJr+iTtS9VPX6vGxrw0b9UgrGkL
h/EjPEHkd048dOami3VMHKNH9k9qzlI0qGPBZ6IjtfJUEWh7c30LWmFfNc+9BLRKwdv0zi/vfvb+
M0Hr9w1VtVBmUsKCTFCxihdP/yCK6QgkRECf7Kd1i5KAmXNJx9zLUBPGEFXvZJ3Eddzl6VTJbe5V
zoyOSNtDUO8n1d2ERSiGzxDvDFYjCo1o2X2f3uAog1B6FbmYyYVyPXJCpL0cucHQ7KUKb2oBCC7L
5WqLFmzLnyOFTSvzCdaPHWCTcQjmhsW/NOdVuS+wsQC59QnJfW/rJtGYjbtXNOpA/olcQCfDvKWE
alLQewt9e14KkHMdyTg84qte4uQD4gRVp0MiKEUK64RYzGni5f+R+eL8fKY5DRAe2l5v4nBSUs4d
qNOY3zOhZTaPZXhuNf3wYeHjpyXTOSmm50ZDp6UPtf00iaj1Hx6KN2qY/krh3iPa8VdBt5ksQA5T
a6VOpFwhUn+tuRhOII14xvtkioHEGpOQ95KF3PITPT2+4f8INhDsoCbT3qALCxlc6LvlIcv4ka0Z
b7iTSx7jeu0U+08zh8BDtYXwh6th2NC0GbpV9e0DAsUANDlzkaAjBYLW6iH9EUk9rSjNB/PO67fk
Q2levBOlJHrNWD7oMh4/xGeadGVJwNUMGurHoeU53Z+VDOBYNF6wDsG+ER7/ZnAWwx8pAKmuYNJI
uQdwF9Tn9oqr5gsbeUVc3OV8LQnr13A0a3eWUAXUhc2nQZubrd3ZAMTrbozLLrt2720P1IhcrhUE
J6xYadU2lnjY/R/i716MRWdGRRe5rCiO69j+Iri3mkN1U7qld0Bd7ONq5A0PDrJ2Gk6Sj6aDSXtn
2c5qz3IKzqNJYRZWyGb+InKGuT5C+8a9bSk+SetInB1TpRU/h2KK35/Hifb6p5m12ZUdwSNpI1QR
BqGpQiuZVc2uRoKNQ4VjTuoH5wAUZ9DDSVYgicXgmtZF2g1/XED1Z4/Rux3el1KgbxidBF3KXcJz
1LKXYvScf76G8mgrd1K2C7SpH/RNufY/xCpcNqgYd4OanjUaOCNdtc9N3nyvmBrExqxqIIac94X3
uSxNgUf/7AU2GKeazZZxwNajMnI+asibhhRQuOmFPhfuhWNV8XM0CuuXk7mo2Yai4lJ+zQs7I9/n
wIWbZQ4jkDHAwh9cvrLSz6RfesLoxU+8UMtZ5aqNfHF8XcQEQXr4JDvlyLHCgeQVTqfvjliFnsGc
uY/7oaOx4pmFDXYhEvM+34+EcqkiubMPhfR5sSbEChvfBPiI4UdptPQpNvXvHJOmbwvqBNpfr4b7
9Ktr6JJNTNNNIk1uG5MftHElIozr3kf5M+QAuVFeiaRflqUcD38BwZv30BLkiKb/hCFjS2jXXK7Y
W3yzZ/E2QRU3iXo3RF/4H19qOJLOFcK9OvgesDsDQ8kUepiwDB8Dp4qe/SY+sHUjeJ0OpPe24DbQ
CGnfsfO3bIF0076ovcCf8HGLnVJQDFHBm0znnHWv8ot+bpCR9uME8OK4jrRSKNWAd3IFv0apMY1K
NlcxmX0WiJODkpCgJMq5poKpMgkNYfOkJb4WSZ/AFTlfyPcfQIy+Iixwm3iUclLbZNzc4awIGxww
UiN0hP1jadCaErgjBbcS009cg1Lnl+gl0OxQ15M6mb5YR5RNo5bH35k5+IIPbHzlLQmHmsfMwO+r
jmgv98oYlW/9i34nZB2FvvbrpVHr7k1LxjD8tb8Bzg1dV0bAYP7vvWUfKTDl+itW2RbtZSMR4ls9
1s+R8mh9BoOYAIYpBp8TiJufOZnGqVry7CnaUFLmWyTg/5CIIwrbnTuKu7sYfW1rC+iB+55sphXK
UqiKDeQ7qmJjm/2x0zgx7odnl0Ld1PqqmDzzPhmlaW1vKd3MpoJ2TimLB989nSN7INJOboM5LQwc
t6odIGQDQ4TO8FnbEZVpijlbHRJui4tDkt6vuf9MH1AbN+tIbjipXFYJWbm+XxMU3KgAgSK39f9W
Z2eRgcDMD7s57wLhgCsykjy59PE0KIT+DEX2ebN4S2Wp/Nf/N8YKgVLEwrGbIjOxmvdj94ORq/Pw
hE5D2FaVVIvek/jTdpgoR9S2mncFZMD31aGnRomn3rKuRpCkQN+uGSf/pwO14UYWZw==
`protect end_protected
