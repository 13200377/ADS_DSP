--library IEEE;
--use IEEE.std_logic_1164.all;
--use IEEE.numeric_std.all;
--
--entity tap_mux is
--	generic(
--		dataWidth: integer := 8;
--		phaseCount: integer;
--		tapCount: integer
--	);
--	port (
--		h_n : in int_arr(0 to phaseCount*tapCount-1)(dataWidth-1 downto 0);
--		sel : in unsigned(dataWidth-1 downto 0); -- between 0 and phaseCount-1
--		p_n : out int_arr(0 to tapCount-1)(dataWidth-1 downto 0)
--	);
--end entity;
--
--architecture tap_multiplexer of tap_mux is
--	
--	--x_n : in int_arr(0 to phaseCount*tapCount-1)(dataWidth-1 downto 0);
--	signal x_bank: int_arr(0 to tapCount-1)(dataWidth-1 downto 0);
--	signal h_bank: int_arr(0 to tapCount-1)(dataWidth-1 downto 0);
--begin
--	gen_outputs:
--	for tap in 0 to tapCount-1 generate
--	begin
--	
--		p_n(tap) <=  h_n(tap*phaseCount + to_integer(sel));
--	end generate;
--end architecture;