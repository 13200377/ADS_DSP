-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
y7742o9/rNyj8Ltbh456Kv2IHnuqkvRWdVwBjyh45sT+78LW0cv2adWsxfNbbgmFJOGkYe8sXZlT
PeqMCNaUn+hROHIzzxGyasPu8z0swB+uPdTWEEmRmsESIWgZCQlEDzkfUxrdBz0JZss3H8R0rcD6
jnOra75/ADZJnIiqLoW51JjhF9gYIWKVvrALgFvlSRwP6Dk/+gHyShM7vZ4+BRMWFTR/8zyaiEOa
wCB/rLUlvSHXeWKA+Wg0/+ARfs5X2eV7meTOHxu54vMFkOG+Gb88vCHbPvBlzoMs6L0rjd4KhMaq
v15/b5tTmkhHamr1+U5yidatTkhD6BRA/2UryA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6512)
`protect data_block
QWb6VSwqzBhbT8yiWaMXu9HudxHfgt5655J1rBZqfhkbKES54c/JGn+FQvEjjxhaPnzMesMy3fZs
pAJSC8LjnpZ4/u2grdyLT7f1Fg6Y+0+nFTnsfcM1PHJiCcLYwdaSFqE8VpO7Z3Ye25NzyWTB/roi
hVLgrDh7/n9lz2fncqIJfO+Nz0xj26TVpCLL9xXstSJ1jiSypRCR/om7g6PCG7R8KTCSGGmWZ5HS
a6nMv+MA4cqXJij8FI8J5KBg0x3x38XZacCo/FReRg5tVouY+rfEEVEecnN7R20hQ2XUeyWz0lgI
5wuMPP9AeyPDau4+OOMXfhL86yUgPilaGn7P9wR9Jciv8KTFxZCOV9CLNPx6y6Jy/dcnHSbHtqSl
ec/gHCZQby+1oXfu+llIR8S/WlP1R1GafV8jjRWl2WdXzdykBO6QjhzW71dUCPB4ak0DwDR9bUlk
sccrBMzvgtC/dL6aYeqiiHhRr8bkK6BqG8tU07xOj5Elkd4/ZimipAIxaeNU544XchEsH8MtmZBw
L/DR0AohXEp2WezLXHKpjSnYxVZxafXTTxUszm35r+PNcYSs2zJWphOQ+uyLulEry9tvl4gEZ/Q0
r5CnoudldrgVrieeOklGgUxYF04m1qQSIDKIa+0qiXWZntUf5munqFzXI60W0qfVXPD8AXT2ikW6
6FREkMslhV+BVRvvZn96gyeCJjb0CzTS/KNKqu4OsB3nsTIrMf1vdSEWzA0zk3abP6urmYdQ1+ql
JhBIBN1AyXiVwz7ntUq+SJgr/uhxZKFOgzrUhJQlZVnIJtB315GA2G+UFuysMlrn/a/id9sYA+03
zexWFbx4rtKWBlkq+gaAzP3o9sdY+HpBvq9dmH/CYcscQfB/tHuUVCqdfveXJIXo3BBBcSrXLHl3
1s79ugj1xBPVXl5yBt5rooY/0D5PM8fKKLrOKjmc3dmwDQpbdKUWuSmWGytUB93QD8BCEkgPLa6X
9Qc+ZuzMFTUnLFjloQi2I1OoNmbsOjecZM8mCH+naTMB31qcqZ5v1W8ertstMzcf6UEk+2SiIqej
4vbs8+AtJgwrNTOhf33JuxvB6QbHU2xcDCovy4wxWBTP0r+crn6BAfUUa0B6qHSJQp74kUMSCTWB
QpEDB+89/IKasr6/YOB8JKtNBlwPSEMjUF4vw+o+YSJIqNO+CT21RjiNxp6/h6R7cWIdfAI8QaX5
HT6aL1q1lYZ0FYnYOVVO7sMvS+fH/8n6Ispal7HZjXV+0DwSRQIp+ag54v6zTuZFQvI9IboC57iu
owWaj966pOJJG+v8icKI1k4gP4LOr2NO/J+8Dm4CZ1yMR0+m0kCYpnNxZhTzb4VWgt+dlSdPkSv4
Dg5LMrWMfqIpj9si0TsQmBhCsbpGYuo2mgY9AZg1wGx1HTturNFM8Eopr4lEY24bEqxctn+ix2F5
Ixhp3TX12b0GL0ENhXhzeJLp9NvpoHJbTSWAHZGdyHw6OBVFjHO1XRV/yw+IDXl2i4VNkOtDwREj
PNA36BoDGwgQUkgD+2K9npZ4rq3vH9RYNQqdBx87D2ZbiuFHO/MqfLw7s8xhlJAkXGU0xzJ/J+mA
az+3Q7IbP6JKKFCLdNMzNHQAG5Ix0KkYHnAXv5CwfC/kJlA44WuQ5TqONWgLYffrgnUHhutw4WRl
y7xnUQ5NRP83EGNMbHjfgNQGmU4bkfPW2ii27SbX1xnqP5QfdxdNUiW67Hr+b3rexB4QDwJgI2sX
rjvbQ/AXXWvDunkAt5WRtMIBPYXrnPLo87K4Yp//6LQjxre9KI57M91hmQqxvzHk/fGWQbsw9x2n
LWMY6kAGs+SMnoGsqYG7CcOiVzqp/CJdFqWL2im33+YF3dGxyHHA8Od8XSnjzmdM0nlMtys4Ovc8
d9piQtnZaH0VvQajBHcMAFFnlF1M8jxtK7txxuUcajMOQg+lLpJJEtUna9Kt5AZwtBgr2ArQ474Z
nYTn7iyetV0YcaV9X8qF2QUcqmNcYoI8aRngAKfhFeEApxOWp4s+y9MX6cyv/S/LY1PLbTh/atgV
dt5LYBvyQrBYaDfeMppS1cjioGKnT1OJnjJgVp6n7f5KWQD3xCHiSfZGejkOOZ9cU+Rx7Y+zLi+g
kLqFTWbixHd7wtl1wKEujO/44Srjlx+TxkwW/3ljroAKNQHtutXsfrVqJRTTMmzmHu8+a2LNROex
a/GMD7fpDK3Jugsf5ZRI4jQRfCaZT03j/pzPsg5kDuP2mGc2ttICbdLsEATCHp82y866c8JmaTgn
dKjKRVRydkwvjVXnS0jIoUaohuyjYGPV1g/3wbD3kpTKnJVVZlPsEvaRlMp1SJqB3JDSNDYCRjwr
QIM+MldSOosKho6JRvXW513WdTz7Clw7e27IDozVaeX+KNnCAQgYzTWHbL1rYaiXyGyOxy/jVQs8
Chl6c0LxYuD50FMQ26hewmxRYWZDTAlNGZ8EA5TFa7GfAgY9QM/iWYXoeJPVg4UMEAusl185oBgs
Jb1TwIE0aEO6R+8oBxTAppstnNeG2JdqY7rL5FDoDd/72REfLaNWaiNJM1fvU1AKNxUQOX1rRhzA
VGoQHfh4SA8xxRYf2wSHfMl6pddd8lRBaqb4aLVfg4/k/zYT8O/RpVe6WXT0RY7L7T6D+dw5uN3N
EkA01Hl4pxAuq5gxyL233RB3XXhACQdYAiRC57LhdkXf+DRYtdd6c01Ws/c3do31Ww4WRusru8sm
btWlpZlQN/wWvShhgSyQeOf0nfignsYBlXSktVgx+DJrKr2PuX9vPSRAMfmHiJvbdNt3nH90+p8e
StyS2lAzxRBxzmMPuyUBjtCws/zC56T00yVyQX5FbkWo5cgE3YE4M9hESWiB7O0nYyFVREO/TVk7
WGFlviGfKegi7SYFkWHis3rbzc0x1QdPSY60bzR5DALXWBGNzmdJ6miK6LHCk8HfTl9MU1XSr+++
O0TdY5jAtY8g/sDnw+sRmivxHw5gAEZJMOxR/jXIVq2fdY4mHJvl1hshaYo11dHrgwORTCK1y6Wt
XsKuLiqQo9mGghJR6hIiO8ZwEf8u85SqwPMs0NIdWDUwG89QiNWs4Rlm4bmdTx9SomVsjVyXPitE
yo2wE1P5bmQb37eFxxMSpCafoPFR6/6BFV8KlXDAAiTHJd0olkThaJMcSkU2d+E0j9n0Jt5gYkYs
fUq5wwdo6Sdg+/uk7zvooUpTlvN9g+UXPw6kGJjtPcwLLlmCXOxN8WgeBBI0tNWtnIcCyW7oNi5e
fqfwoOI2oPXIP2qu8vRTg/C0TdRBJo1lzM348BcpbqlRD8Wudyd+Hu+OCPNgF0ldhI131ji8N0I5
mdRI1A0z8FJX2B9URe97Iu04fqHQ2zpIH8IKCpvZ9inhVwU+H+RBP7fW1jMtWCOBPuuaPVIHmRqd
mRmsNq2tF8qMHVAQGdyfuq0vjLENgoLz+65Bx44e12sHDBZfEBlDrw7qR0vUHQ87tANXYpuR/0xW
FDbEV46HSP+UUfVyvT9hXITPeZjtUp9b0bPUUcCXtzkJM4+3pa9ZZyL33/jADtywDHsHegD0T0gx
9MZV3tTq3tDJEI1WzMt4a6b1tkc9+d7EW9+3FI5wATh+0lmmFauh2VA+vNhx3F2asiStCeMPGpdu
RBi6BEqVBg2Lt3uZMpX0QO0W9MQUtIXfluNAjmn+j1n10ZiLccAiWuweOS3/93T48R9BIllA6tRQ
b8hh10Y/zLe103n7H/qh9zxTzXIs3VU/P7ENi9oX19fSsFqj2BYcq0OjqfNOjj1q5vACx8sEkXqu
krAvppy0MFnv/BYPcQ+/IOK7TWsO8K14rQ6pKeurcuD9q9QvdTP3uhm7kBohLb8Mrua/6gPk81z0
oUKnNmLDgMfnX00wxesOxRUJqJM7nyupjJaXtdQndIfTdf13fAmiVsMUIesBSMejQihfKSMPjCTX
Z5Ap5ECjsk8ySSimm3l0IUFLbV7KfCLb9s/4uAYZbmdG91DCbYz03mEtffnHPI7RLXBFLDeiz8fU
O9twcDhjvKK5oRwJsoDfnWAeTNuwrK4I4BSgMJWiICDCwGVFgLGfLNn8r9Zow0bvyQ37mdD8waFp
gMmLo3KCyTnW1yB3/92HyQ+SUaEiA5OcITYWal0j290ZNIzb0s+lCSmDMHXIJa7BqvZnVYGfsWb5
T3G9rBXSvQ0L8xcthp2wR4SNFyeYgU4EzXF4ULpsH1g2I1N+atPEIm/brrBF+DhlZiawbYetnaP3
iUBRNhP6X5VqLuQ3nnzXDP8CA3OK8CCpZqKT3LjUOpGioZBXjb5Yix5UPAYqfYIW6WTaO4iXHwoY
GF2EeZS0USLDo6qLrSCjRtjaFj2t0a8ZzkeKnn7OXnz3yen4qGr/rRDRlQzegMp/K6UOppz6yGwL
dcX7Uqj1zQNShMqFUf0LeCgrbelNmWVs2DHMGTl/4nGRpaH119v6NBOXEX1e2bXw4P+RtpOZscZ0
mkEmvqCrbRAqSYZCZc9a2lnbxqLUWGzhFxsBwwpgztjsBa3mM7camsrpYlIqDY8z4wJZ9Rh5gbRR
ecMcZ96R6A3ffhQJhiI75h/iWmUWvW9aqDt7UL1PRU5+ND603hWMNZBe9BKF0XmT//Y+3ja16cq5
Ntlpk8w8GMXwmROxj+rWMAXt6SUc6i/FsbtS7Z4pT7Tq/9ZZD5Py0BozI93t2G62E5OZ8B/no1Lm
v+GFg8Dk21aJT0pbX0nvqVZgvO8BNoVVc2VuKAvolr5kpLtkmBmOEeLlO4A9GHEirXzotOL0hj6N
1/MfBMKf4iwedxei0zMVNZjynIosG+95DdyfzEA37z1MF0UeswTFWLZ4byI5nOWQJar4lZKTr8hL
vpE8deHeN2egnq/O0oDwpHOx1qhX1rLwnAfPzGJchOPbvjdF3XCT8Z/um6YHz0IYNikKcOrVRgP3
YkySAA/7pDavWQAa4CsjWwRaCw2V0N1W8hbPT1EaUzmFPt0anCZzk084vBDEMUsOHmUsnJphhpNn
HLBv/lAk9TUsOMstLUKvNpoyOT2PnFiTUpoLiYgSVQ1NpwbEsn1uex4cBT5KN2uTJxhP1AfSX6Qz
r2V0zL3SmFFPoB4ruYlE5qmP41kwbwPbKjja1gdeHKCH16XGtJ7dsLlL2BRISEbgCQsF1Wclsb0I
vbIXhs6wi70tsNv8g6EYZj8dk1jrrJ0CBgPmwrvepqrrxuCucYKf/6/Sw+Fe9b2PBRe8NytcCmfc
Wbfs0XYOktbbQyzmfe3K1I7aSJiUHEiH03cO2hA+uudT+MhnupGDayvJ/Eo8qATvbYgc0OqiONI6
gDiNAu0CRYn5NQOHI+/DIDyRlVwQoEa9mhpLeo6mwfzYMYjKhUR1FfO9VnuUe/kd1rFd4G69Cq1t
OAvOmQxY+xky/ftpV0XcU1T3TC3bA8g1EmRYRqWi+iiLXQyBa2gAGct8LlWsPe4W2+aQssvGhph2
5xOQB9Rs85nooqfg6Ja/Uy2/ZnExMU6Ct/BSQr3HmrnRbSgfwDvQ0ghGhHJW5+C6hObZXkiPTumR
NfCoJ3TzMH1fAPQcA5LSTkCZjdM4OdifUDrIE/LOY75RMM6/pOwPDVFWhN+lpsjDmrcINj1Hi32R
HXt9H6XBL34yDAR2e8/2U/Ox2F6G36B2hLw/EhI3Aig1hiN0V5QU+i42zpOGoW+ls6vF+quNGG16
o9GNNpVOT3uwVkQoNKxLvVd8OwLnv2Z0YRAmM/510h38YDOX0Vh/L+1rPEsL/Eju2fRPRDlzGSy+
Ij5lWy3y/wWqSVmlq/FubbGhkO/tJOa4Ju/4bTaM7SVP+9xf5Wz3HwdGKt7yND/a5UcTFHZ7QoNc
eboAYPuTvBxOsBs2tqQ5iEPndC/nWkxjH3fjJ7qbgHAyLJXnnC9KIYlPA2DwY/DNBNmUUp8TfRoG
hE+RLPsNydyn59zAxwqXq2rnvkZ1+nyVS+Nor6DwRciu2KagUHzbL6epHpJNGa3i+TUVawve67vg
UeuXkyFKs+F+YTHXgenVcyJEyzp5bLZ7h0n5I8cU5GiRIh2wdeK7NAXzMU6gNnxDV0+MMQmcyDAa
kAgf5OvZBAkjW6Dkc/bh6ebY4QfeJDeKoTXF4y42FM4NtRO9P4dXc/n3SxXbunQurXxwRf4yyQks
al8rYYWmjAf9gn7ExWoDLYwtGs3gxXR+oKkJYwwGeDzZBCYA6lwNxpqFj7sedmQgmCotwKEBRW+y
ivEWhUXPgcCtRoVDegBp71/0/e82Oq17n1XIfnO9K25zts3f6t/frh5Mf7YlSgK93aPGZAVoLpwz
izsCytS2mqLA/zIdnRbspBqpIWEq9apEVlMFPmE/ueCx7HQSoFiJvK00FtpIsum4N88Fzw4nDl/F
U6iP1xoLN9XonQ1iZIndana08dLTegDQ6LJchawGbr8yO7mYpA8HOe2gq9TRWNRanEijx6cO3nMT
763EQXqZGoUbX5NGh9ZZZTh35dQkUloU3b2sjls9wrVgH67VXDvEHEZcDqpFN2Sr3JTpPB6bVQ9x
6WgQ8MVntLVi3N1n1JSkK5Fxp+Rjkhvdr8WiqQhM1Q9zzqbs/CVrnKU0XHre1Baltya7K/VeX+oi
BzAelsgZ2agZ++T2ZTeH04Nq3p6GgAYcbAInZLxm2PVbK8NedOZnltqwRFVyoFev74oXZ6XZPAHT
X0yIuRbncKicLs9j9vRrTgL0ySvChPpfw6HvYA1WZttKPjdaZ9JhdABziS3cvzt5hotp0R2iF862
YJv9soyZbnb/JdMmBexHkzJ+Mj7JfDnJkGpnanmkMV8il1jdGNzEEP15Z6P1WJ7gXAQMcjrTxa0l
AHzZVmyOE5i5XLYfXIN3oggGeTyFBQjiJ6yCajp2Y+5xV9CE+zBi5Q3XaKnTEvh9zVf1QAgtcNb8
/UwFWKTiCPHks/60B1DX5cqeqcADNGuyv6ELsRo09owic03qnfU0j0CVrGi3grREXg1mFIT2X9XG
2imtR+yH5XM8JfNa4VaO+XaUP+leODVCI9xzHuHJSglbqTaGLU0htGJ6NCXfFiUv0FjwMambnpMG
eZub6fPYbQVtfikglGTRlmkwXmjvszcq+FDWRs2m7LSomi0xCmihLV0SmMSVx/m3j2/Y1gOXDWwq
cVN867qFCLzXJkeLa4ggqXpZbvZ0PYewIKnqJt08ZrDq3Dr2uayi6svC96ONOrNwL/d+Nxn3YKUy
B30C11+txN2I3+tW/aLMR1D/GU3D9ohobfdObHBRXyKZUMeK7ACAr5E2bNiKJMcDZIEefKqAMYEu
vKDvfDmV42jYaAsqx0+PtdeC2vlEng2dh83lI9XdMLSbMV+tnuAKFzAauoUPXQbPd9/4bs6UjQCs
oqyb4fz4WdBU6NpHGhi7xWWxyJqlKffAhSYdnP3ePQ1VCdH0UkHos3GOGVkGqNgx7aHLMWlEaT44
gaWxSJEzVa+KS8YAsezvBjjkjpvYHVO5cY6lFj9Js+Msy+ycvaXcNvmsDgeXgZuKc/JkH0GrLWjQ
FkJmqF8xIQtUv0UOTacMRA6zxgSb9DCjo+No7thw8UActbEuWVe/ZXrKWcjEwDlRpe8/cc7mn6O9
zONVg577ZzfJaJZvDcgkm8kvxMxqMgaHqr2SMi2+PQA+jzNjONFdAtoQZDosU5aHlGw2ydhT2MQD
exavQyLeBOQLs5cQQR0aSbeYDBfqF3GzGeYxgIAh2xKtAASpF9LPrNLWLMpopIS2YTb+gS/wheGV
AlpxRf9vPn3cvBzi0n5r9cwDiEf3+32YRjeJOFGqs8AyEcU1pQHSAKGB9bIGqz8riQz5Dlw3Ix9Z
DpABaiohtSPvgNHAV7bZQPlHCegpbDghXzWSkG0NsK+q51amCKFxEs5KWvbVelZzyP9tkcNPKP+Q
pNh2jrsRQG2d9INTTcRHpxhuOyev+e5ih7ui2V5YS7XPqPqUXWdDpQimnVnjY9fj2LgTkdd7+QVY
BR9ieZLjafGMpageubInYtUVwL7gmfvuiVHKGasH4JaF1CTwzS6VNh411yK1szQCBaBh6H9Zlh6k
lFudduQTMpv26MzcgPztHNfsoZaCcYimJbq7K2rBD4trmofvkejLa5SN+W77Qpre5a3xqCciTeT3
DZVcY+i58v4sB+jFadP/NWOaucZyuPil9eJGB7d0xDv1g3uhV21/U+tvWcEC6B9Z1opGvuNrWxrN
XrxHFjVUypmaLHnYG4VfSV+9RCXzVO4vy8aAZEslispBOYsuKGZJwqaBU8lRZfiiFVjsHftlqgfG
OMX8a0+u3yo6Rna89zn4QfA35hc0MnMOOc1u6cnqj6oxaenL+7GvCb3G60CVUyOZBZwuHbwclXAI
uI2EjTL+W2D5enwYsxoGn/pJDUmojkEtqah6JobXDO1ww0gAv1zzSoe7iyfArzQ5Cqjy7Mt9r8JM
pa4YdTVXk9z2vQ/ZuFqDWXA0UnTR0aj/RWw5RFlUr743EtdBaISQSPTXz/+M/iyXmLtmh9sXaUaA
mxEuBq58i/4QgxKjBoyZP0LZfK/kr0tXb8yQZ+kpW75fsjYRVQFrD1I95VyalJSHKjVwt7dBVQTT
g2CDWYYscpGDbmIT9rYX0HvVMZfTjtvM5l9xvvHQhW86dpUiECYJhfORH33cD48OZz4efl9b+IH5
ZmzjtbbkPc/q+O00rT0=
`protect end_protected
