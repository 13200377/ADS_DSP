-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
z5CbYR1nKrdMSOJxi8+vgJSQjNrdb5uIddilxhcmVy65GJI5xAXvL9aWKYNRcoqh5nN14WQKomcz
I+izoleuCR11JB6AJ6X/Ha1/Qfe2nCzXrbEbNoir254ed2F5pe/EdvKd5Axh+erEQ0ztiYGy0x35
yhUF0bJjHgkVTtWMX1uDrSnuD8NbFU4Tz6to49041aCfacMiVEPrVPumg4yn20y2DCN9KfJE5XW9
e+XFNGxJLHhB9U3QNK5SjpFKEpV1Hp8Y8xXIi0wFkjJXTcp03OqK6mNGOpUB7MFPT9/knUH+ECEd
UsTIMcXvdegLVmlSKfwkzCf+fx7SE51jX4FVfw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8208)
`protect data_block
B5U3sSYkR8Imsio6/D6AqElzK2oUXrnd2tpEZrbQ77pscVFhiUnmMMZdqTi4eiTwmdzs0rZP8nYD
X1fetRNVsMtbB5tRny2ERRl90iIF0MG2WiSQ1+obz3KUo/KrEP8ichListvj2KeHKVpVeh0ZlX89
EHroZnj5n8bN8btY99KObHjHPKVw7wI1LWvrDZCny2ZXKOP29tea6KWFRaOB2N2ppV9osbTzFQqT
pTP8CZOBFcd7Rcw5w+xMXJyXG86ViHUCxDSUQrgdgQBuUc4xlru/3fw1+oKBCPLnRYJu+iQPLltE
ejgSN6084ArWKOiqyW9SAppHblzQ/KxdKPakzms3X3OhKtAlZ+EFwCH4R0YiGpudN3KGRTUX9p5n
Qtd6DQHX8W0xjXBPRygiLM2uBamvKx4es8cIzMKrcHrek8kRuqsI49+tCg+lZhT8+BmXhGgyQXmk
RMzDa8XKVqlBvVUfMrVu6zFMPgwVaPDR4+u4Rb6T7RuDB6DfA0EZdIJ2sGHsO6HjPlmFtCVjHS8H
JTqN2/FlTdSLYYx4LBCYovjguGDeFwx/bnJf3et81rJdsRpt4zFPWqPq8kWIwkGTm67rWUD87DoB
yaBhsd2SBAQQh0Yb7V9bJz85fQqsvap4wlYO6AVzG68ScjMx09B2z9ixhA/Kpr6BSIt/pOb766fK
5VQYPE86j0S8yh+LPBQkVMW2f+IHGzUjSE14Z5VrqQOIP6Lccjy5Uu3IwUnm8DFpwnqrvzcTpWR+
atwDNJFO5IHYAxjjJUDyRGSoZNluaot6XdcwiSxvAaoi/I6cSJZdTc20EdzZxanlwDHosqETtwtU
yLRDrBFBZ+6HRf+ZIGvSt/3rrKg+LTgraak+DH8kYzAfLGm2glNvewzMFuaavddEMzyK68u2wlyC
2tHAco7XcWQUFM5F1f+O/whhpu93Znm4qfVo5/dXY/Mdyxf5DjcsNVD05FfyIBcQEhzkCMADPAmg
bapXLv5oIE5OyB44pc5X/EiA5Zdo9C9K37TI429Q/9kWlF35t+W/P7apgl+7EIJOKmJR3PLcMbS/
SNknrj+1i7kmbnZC1cmMYtV5N6XiNCu695Dh01zfy4ePwA6xvj/lPZDccu3wBsFH8xkY7tLEVgcM
6A4iB1iWuXmz1+6huvxl4S+p+8ZIojjpqjX5CPHJDzQ7Wx6oEdzqnJpKEAS5U2Ql9hqpfPSXs2EA
NHfESmYEBa1m/wNvyuwd1K1rgzi4GeY67f6Yq/xYUwvkvzWs/7YvInV02N+QbHKA6Y1zQMforXBo
9iNeO2qbNJgdGDhqdIt2CD3V1NNyPecUreNP0MSMucF0Kw/HO1PL6hqWFBuS2Kn+TW7EBaccgTj2
9KLrRt5XmLsPGo62yzAkOrQlVGozrMNZD8qwLsXcuKW7NvW6InzUGjNqm0B0fFYtBb6Kmv7cJymX
kihIZqVoFrxB2HDCb4YayojgivWtr110YEnxTMRqvdidFwQt3jontOfNXQYnjaaIeV4rcNMaDCyn
DmR7pwHVDTbjd6NSwj+6VwjtbDf6pkGno/LwDvUzulvsloxz/QgnS0zGW7NmN3t4c0CZoqUU/po4
0rvCHduMCn+J1DEhCJwJlNq1FH6tEASW1phNA+ZAQ/+tPmMiJmGCyhZjh4mXmgO4NZ/pQUUCVyvx
Os+3lWnKFo7yeFQmsmQHSF30mPr4vPRMmmO2rxyiq/dsCK0CFzp/LgwY2/ksU7egz+ls+8vR8TdH
macKwtyZ+Nh+rs/oPPCiQunM8WpJGFVwUs3f9V1ysmCz2/qwPeuB95c8gP0RgyuJDgFRjqEkGRVP
+YzxJG3utVzWcki/f2DmVEqdmZE/6OWmom2tqjxOjElQiFRX6LLycv3mYEnj/ml8hfx3YSve+FGS
cSCOg+9RKtoaCI3u0wu7HneFR7LbqTItD6HQqFKHR8il29ND0PQvopOgeqe+gP96pumS6iMOm8Xf
spCshbsWOEdRdN06MP4GxLq30J1adSvfgyMuzAOKVeYbIaX+fdbGJ0phjBfqoyiV4fY7Q1VOAHjG
abm48jO1rZoOCKIgiJ91EKwuAXMtPnUt25SilHpNF5qaZxqlhCNL++SmkSJv2V24H7kO5gKqzVTH
liaaFr6FcdihjeKf3cUllYZ/SGoDFz6zbfjBrNgKQ39Ah6tKMBqCC4k+DonkA7GHxunys6Hdw8vj
57U3oo8aogtWIV9HuFSgBnfbrFg9xYLbNGY8uepnoIQzMW5hnfy9Uo8SEuSZvfgmi8Q7vp8Yj3KV
6AIKlNqzFpog0kBXkBaiTpIuIvKZ5k/l+pURxtL8MhhTrMIA6hFSVLSmdFmbhehaeqXgpe8L2qqR
uhC9QuYxZdokslLhPAk4s2AiE17llbPHTWACX4erobkrwps0JvRhjuAVNDR4+rH5txkwGFV/+VV6
woE3+qZMgi1WkB5y8lxbseuJhM/FKKlFEwe1ye4s6xOe8AvNQ+0EhU7CJpU1HMImJ6ty6p24PVKC
dtGE/w35UQi9HKP0urovjmqju38FHnAhy0y5Vc5y1qSQpVXg+gijiinh67ynGrex3Hjcawu7sJR2
sYkVlX5zMjb6mdwCpbQhkR5S5gXjlKB4F76+az5bljl7PFaQsnpPaa3R+IRVQvjlGN4T9wqAwP4f
iwV0onvZLRRdmYtu7FVI0LdPeRhGZ6q4dvt5J7dQW+dsUyvf/kEGuNt8RV6LLCpTEBWU3q5PbqwN
XW7UrQs9CDeac3FBA2KFx6hDJVMLV7jNvB7MB7n2U40h1h5wgSHqVlykiTmGmGlVmnnzDwdXQzuA
v6zz7Ho/F5ARKG0o6bc/GhWmVOmMO7r2lnZm1vqYtjxGSp8GIW9FEdNZ3JyQs7GXFN4tzha2uR7Q
rbJP5Lz06prCdrtK6lJnN7GsUwugzORqLHikuA8u23bTvzKjjWnXJZMDEY/VZPcSyuCzjWV3pR4K
VavnubO+7jMcGYnhPDJ+Ri3sexVfrXU2wmZPbypLUd8xqghRG0wEKOuozQC11NMMwS4s8YRZrYHs
fpmaguQNwvAwX1wYXkMFPM+ateXz7DDKpce6ghmYMrvolPnNGvhc3rWrpvWIzIYXLN7tUdssph2r
1AJhR+V1VPOHdN7KF1W5giVKom+V6hRmalZa5xAAnf5L3B95ujQC09ujS9GFR3CRS9eUq5+FAJJw
j8iKr5lp+8ZgmRnku4s99lAqdaYM0fKs1EGQYUAf2BRIdQ95kNt5Dlh935lGw5V8WWVSUFRs3maE
tGRchD4mpXvLP/Bmh2rhhC4oxbwA90irLKuij9LzYwT+3ZhnhCgZhqnQWE1pkn/P9VEfWHoxXzM7
Vf/8BKkfsFiJZegcZJfVRCCA1s8wVQ6OLWX5wdedlmIRNHlllnNxakdUIzpw/9TApofz2XgTUT2/
Uo4BAPN6ylqA+NQZrUmI0Cl0a+2gJRbxExpMBqURl2GYmNM0KJxIN2oA0Fhz9OKZ9M0UYXSW2Wng
0uVeBUWHtxKq+ZEUCyfHzIpymdNB3WRbDvnPlz6qxoL14pFd0BVwHn3olKunAAF3okEJrF5Q0iwS
Ky7VtEpsdde+0T2CMORp6G4ax4yiCTaCr2ULkj63FDRx48fS1K4ymI6mbljI73e/5LcvfaLfzGiX
1HJujGq/w78OqpxGtvWh8LbWkjJ3rYGmu0+j53y+IcJYKOzqofTiyNVYicYCYAaS3nHTWbR//s6+
Fv70YnNyAi36L1ZgT3iMkssgZAi4NjYXi++3r6JPmVPtzSfBN323IkcacVIqcppF5oOGJjglJlPx
zXRJ6BC1r7FWbVUdjV4RZ3kuo5lEJt7+Eta76zPiQVvQ1SsoysUoqOIisscQ6uztQvZp32HJDIFP
tk6pS6p5a6z5n+v9kVn9b6XgBd7FZfz9XxAPde++A0CRzJ5yR9Qd12Y+cT+u8zslXA7/UVO8FGg3
nifja/o9ozH8QtGCTlu8mNtN0mmqDHnW+Fr+IShwWjEiEb4yPIgNCPUMCOdXFjwQMzOBzW0oZ7kS
lGF7GPq/fjIg1DBGstYYGIVnq/uv3E5EAATdod33fLn2lkMSnSp4x0NBbsu6CefzyyU2Vkl9oPgr
YLP+WO4vKy00pNwdv6zajPEiw2KxSH3JoswIY1LCkmZD4YXQQ/ML5BjP6PbsCLTc15i4mvOPmg6a
033J3MrjAsheq27dTdPdH12ae2pYLQFvH5VYaRY7bDnpal69K0cDE8xjF48cgT/jHsx/RIWzRpj8
S+KADhhUd6TWMBnrgvsIK45Xpqh6nnDkn/oKq8aTNuDurs1GPKT+mzE3i679+ZKMUxCCil7zbbp3
0MqvvCZ1t8xX7YaU5zWGJuCmCJmE2jcZ573GOXBoKNIxbOqUkEQyjz0TIuvnlgbMXNE/l0ROoYWQ
JUPILDuXj/mU0BLiZrKenoMlYOPZ+r6sVSnlWEChQKrK2DNpv4po22zdhirYDsyGxdrJOKCfdX2z
19513DNsA5iHHS+38SrBSz9DeCnrA1DpXJm/fE0wbtHn+KyPCBSl3Vzcwqp+QnbZqDqI2bwWW2g9
6etvDpR5yDRBO9sac7Xw2kJjo3H14WMWWQbRUsTMOQwBwcN17sABSi1x9XGetnzy8JjI2pyjweMo
rXzg8jKBo+SlS9jpPxCHzjnho8ztnqzWzwDZWsLA5T/UpQZMu16mqgpOEDIPt5dau1UviW9CW2GQ
KaJLslxcbCXFesWQI6fuutXzZW8oCgRHVdw4ew2BqEij89hRzZ8oxphLGTbIXmrX5h12pxobM+Bz
d2OI78nHWfYy+aXEDC29g0nJybaFkhibgkrQPiN1GRtPmkx9bRUb3yMrmhlNhBVTxmAtjBgG5xOL
NFto/5e1jqkgs/kFwaH9MPHEJMP9AIghZn7kjxNmqsih4n7dkNrYGKdgiL+nlffn5RIud55/vpn+
P2OrVvM6JrZ6Bh0UUMIDFTOEe6SpVI/ieKj+rkggC+NdYPogSPTNEqw3tNFq8rzrouuPicsday0P
w/ZvPlXkz7JTJL5YmOVAhlZ0e3bUHdbtvgvX+fSP0Z5CHXBZEtjQXHxX20mgoX2mFpD3gbX/rWTP
/QX5yCEuYcR2VfSuawwoCw1AeHg8fwqi7EImVpIWmUvZ5s77fr0jgzkJodwyDhfk9nhr+b968SMT
pJMN2fjjlojZ9bz2D0NMlrlHM9ng8dv7ErgFS/1Z28t/BtiDtue0gqt3Af6MGWoSBPLZrmWzz9LL
bwDcCPEZdYZ91HGI5EMX5tISOvqrUekPx+ydTULZj2ySauRnb8u1KikqyB5rHW8QjHEFp5vZjY46
5Qou1yiaQtaAJk/Yco5vWuBJuYH6xaH7RM9UnBgLplo3zcOVe1/r+DQ++bjcfuJDea3BJ7OMEwiJ
5b0Dbnrp7l4XWMmuIiM8Jv1n+IAbS2MegZxCIEUEkxEuOx7DD3pFZIUGU8NnbkRFKeWsCnSsD3xx
ZkRejX+HrU8HayQJNTG4mY/r8NtM55NLWIMkGth4XqtKZynUzUf5xzLMy/X7B3ppMU/oPg0YzgtQ
3USqhnM8i71r5IItm4Cm+DsVxfWWF657z8acw9JQ52tygp/MVRyp36c46RUs5znov31pKpjRCXZy
0Znmkw8cXqwP8Y2irj1OzNpjgnR2IVlOeh/1US1bENY0QDahVs2YLTl5RJm/v/kFpKAxrwPkO+ML
ziRBOhokqFz5uci+HCKracvjQkbPYAYJ5TZ9uyEt1Fizmzq+HN2ZzQvhUnbx+l4tiqtoov3i+Vf3
GCznaGc/Qlce1iZtuW6bPL8mk2TDlfHnu9Cml6cT1QUang0gVTGDkiBwc+ULOb7xBgeqovFSc9Wo
qBEQ2klmvQakHur2Yw/TEf+ANqBemFZyMyXbTEoSDquVGPEdL6ytPHZibaZdyhx1UJ00M+lgB7OC
9WSBKn84YKtjCQzSz22RJlnljegJEGJwbZm4BVwWFBGe+BpCUasDuxr3DyssSEz9V5Of6/Gih3Tf
/+4pF+Zj5XG6QMRQr5knMav3QMpV222ohohthb/64m2CDAyuWVcJNaWYevDCPSZek+g8klhtY3yf
Qc6FqmSDgSKtyCLqtAV1/Hja+Xc/IvOtskFM/Q5/Oem5P2VhPnzlSYyxSgm9Wllda2WlRMJntReK
Ha3jZZcJnPS8l5XuCbK54kxKfhVchHAEJLqh2RtvFUGCBeGetNfeu7mMVyYX1Quwo+7RGI/kEO2b
hKcvsA5FiGY9p9Nfc4YGXiY1zpfm7WqOr0k7OJI5bWkp37OM/OWRHxU1r5zX5W4fyBTG5Or6yf65
Djz4xwT800cqHABnFG29Phke88qNUh990+yPXT/PFPG6ahrvklyFioANkWa3AP453JIF1G7QI8ob
IYGDR68MkPzvZApQQgFektzMNTKcx1xoiO1YwQmbXfoFq3AEl/oDZCDAXmku4QqLbWA79G02yPLY
hIaJvyv8taZOaABU6vBVy1yR+tSGJ7dxe/dS4iPw65BFe04GDyZ5KWu2duLpGXR2VvpB56o4p0A7
/zbe54hiO8NoVD9kEW5VE1b2BIeHqtC8pI5KzzVOXQvc0THrvDpqXpnjB4SPZG2kHTVcaPLM9c+A
JrURH4wpqdcPy8ZqS6ZNJQyNe5/hOBSmD3eztjKxHefF74ax1V2WWAugse9KEUtFRQgO7o743P63
A0CabX9Y1SHdatrYBzDOATae+vTGduK5X8Is3rGsppRs5G5cnnGlaAqFrSf5M9Ef6wfcXLzvLHoD
sbTGnhW95iGFRAGglOBGOe+BR7Sgls7XMg4jtQ2Ao++h1BNg6mExOtTxiVinuURDhWRs2BPnxiCy
pdftZamK3x3dNdHs/GAtEWeebnfumQPNn2iq8F5QHlFvLyHAKThkx7kS1QKLaPdwwcte5slWIFAK
WY01g6yUexu/fHrAPqK/ZcqzucGlk5v2wqtjgCTyJpQVLV3ZEZeTLWildWsqfLn6mlJClK9X8N4X
xy6IvydxYi8UxuEJG2evqX9t75p4tvjyH4CvbH10SpqGSnYXuIKTIl0QtbqtnYzpQP/PHs/kzSzu
rj56lnAnaqiT52/Ru+8qEEBGkRIYC728/cQyb12ZzlwsC4ZvZ8q59w+SnGBACW37GglFXamlXwGv
VjVeq+dUJasCrwZ/DU+lJfr3C0cuALCGL4Hu3eNtc4S5BT1LO2a/7KyS7IHJ8vWKCdQCfjuPv006
hH+l8QYO9YH+EUVIpi/9CGlm+1Kf4Fsn5vzCMQJ6rs+ij3yBFhqUoIsruX73C8wv25vcbKBndyus
M/O3Hj2XY/j4iK5kli/H+rhA0BPRow6SL7uuAXzR9nN9Ti9gT6LgFytbbBnpwlGkWtNpAQUDb5zI
n3PZiv61ut82M2yB4U23l8s3z3j7SUNrxu7Q1Lz6XZpoG0PiC5BgxxTFw2Cj0Z4ov1Ww4x770WRl
OxBRzH6PVY3/tf6ogSAK8AUPGGLpDcJi4K6kgdWZ067c8dETxSLLwLrE42NGDx7wJJjt+TiJyvoz
SAsF1vu7HGLp4iToHN2DRUvsqECd28OhXyKMeNYda80aEI4kwMuW4oX5Rc5Dryf91n+ZNUmU2RBC
qWK4lRGbdtmA8MbmzvGUEtypgTqz3nuclFnpZHVlHpLEaTKKO6kV7oZitdTCQ4Y9c1Y63+qr+Cu/
BHKjDPHEQaeqW05hFvu/3DjeIMTQQhPo0FTlBkIUIPwSt6sgbyLiXnR/noOl0noxCEgCS3d2BTq7
vPvbO0R+wSlnm7X7tQwXjN4giOmtgxMCViq9sNyK19YaxbKos74sKpQO64q0gGorMugDyCAlF9E8
DZvWtQoIY0vInw3vIz2hwTpYGDblJjXmnrKfynVGhWPi8nRTfjiLJPNItWIZM27wU3k4znzoThmI
FpMgeh0Ube7HSi+md4teZxjJmn3cPDgUOTk47sWIkBjbetppWpnm8ekNQKTWgXtmz32g6J63Ifqm
ITe88r9LlzvhyEquE8oIZy3re4f11c/TadvKs/hJWBngROz1K+wQILE9Uj+85QxE3Csjy/ncQ1DG
TvI9PVQeWPQEToM233rV54M2ey3xeBZpsqsyuDAV3p86WV1B9Grm5nIoCIFfrd6pwEgrBPjukgLN
cv9nCpqdQ7xcOGMl0VfLMGroiI4ngzbUxrV2g+aAGAhmEIypGvpvkzvW+XrKlZixkwXxpTYelUrN
u8xZ7oAqM6AclgPxYhrfl9iBsxPlS4EteReFSVuL8wh7Ht2KzmyEE1e0zoWRFBliEDLCYOlE1Dqb
zUUPgflreh0lrFsFrf49IwBM6d3R6Ovc6ipWlvYjuaXbQFWi2LHfmFnV4XkIvFD6iI5ehXq7rU4B
hU5/ngWSiFQT5MDbp0PkjJlybiLxTrDh998J4+vubauER7tybebCyb4ez8EGZFEoUG+Pw/KaIeFn
pU0BF5TycsGOJqXBxK8/8cQ7OzEVVgp5oZuKYd8vKDU6CnLTDta1krJ2KIbsY8zM0VWJbx6Edw6C
IiptKO/U0tt7kLqmh3Zo8VaYio2tAb8ddHbRCFqpMtvxaNc7fVtP3gCZd0eI2jB9F8WefE+u1wFm
eqDbWWcLsd2oOcz5vu4sfchu254JTwmGoU+DnTWsRg9+APmXGlTU30wPOGi40XSo2qofxwLm6U2M
dBOzzfscQIO2K9I3ySJut+3xGzWuFvYP1OiBqqCM140djhoNslhnz1vM2iQRLHdXBpvSk8vli3aa
3bjx1BbEDVBpEUXXtFGJdCWS/ywuXICuoc4qFzXSrY3lqGUESXTTkn2CSDkFYqACX9QaGDBsPUEX
pM2GeUV14IHnoREOx/G8pvnNVcVIFhjobT6C+IBB1sX/VELvdSvPGfa9MZoH1GfUn9QGnwf7y8ER
1BF6/bZVGICSpJ3vC0/tLFPhzAQN35YGEkYUrHTFccvse/4JZPlQ2lZ4nP6bsikfXHDlgkiaRdXe
mrQiHBu/LKlek68AZRZxSUN/F+wziX+cfr7LKYFK3vT2OCaPEolR1RnnxWQ8cRIM9Kl2bD5NFTQy
0zj9wBdHOG3+WQu4R7xEHt+YPwUAoLJvXZ8FNdELxveRS4bx4op0aHx++GuRfII28hBhCBggbKlg
UgVUeXOEFjvZqyGuumHZEoxs24BjTY2jRKxsHdtkKQ9CHX5l7ocixCXZSvS+5R+jM9/Fml/PGBCg
z4M75wl9zKd9P3pZmxZVtBGbpnn8Ubzkgx7gvD2VnT+zhpNrBIlyKPH7xs48wi17r2DlnHAWQDGN
xdpfZ3D+xvcJ3HzDl93KLwiAkYA+gHNmDpmdOA22u40z94bT/irZ7wKLwMHx5mJAomQa5g2+KOrz
FDhHtQ5Q/9BpNQ5jjiSvXKolROslI9Vf4tfFItpgkQKEMJAsMM3SgSGFlgL8deNeMTXnW7Zi/ogl
2FnHhFLfFy8AQ6t0MWmkVcxjJHEjxegAr6JX6KfygHyrO9wOaCDU2XcBzIdZ9MHICPjicB3mdlYi
W5ZqSj1RPkTEcv3kxBxf+ybKqYRjVmdlrO+zdTSHeWbD5YG6r2cgTQx7mpyAzu+tdQM68SVcPeIn
NsatDuxYaAK00+xPT+YRclujSLyb0sIuWEI/+G5wbaO86B8DRcA78wENquzxl4J8Anps3lfqpTTO
Uuka5RkbieiD5SSc7EFo2rmnyBaehDpYoOQcnkBcoVXJSVnz2ktBg1542iKAEHIGdNPbDlkP3QfB
jp5T90Z9I09CdHai+2AztkJjJVCrEYyFdagY8EnrU4xKLfV1dDR7nKG27qc+tKkY89ujqf42d0qL
FlSjpF4WEeJFt8HZotSuQ8wt4dQtqMFh2irBUSQ3oVW+KI8X3PD2MaBF0O5eWZosIMi2/Z4cpU+m
6bcrRDBHI0gIUNL9kdhbkFBM0V3MpDKn9yWKh7qv39LZT3B5mcDn0nXhQ8MeKQTfjbbrWA2mjbwg
4abepAAdw3ewpa06B++YxyOK3I1E0pD/rPfYFm6ID0cUYOOc3EEtcmPe24h0Iup7rrPLiJLhWTjj
ihDIy/VnpYXGYea9rypNEQY4wK81QnD4E2DhEFsFK/z2Pcu76P+fkvOMPjteU0R8MEmtQFTIGeUW
xGFtrdQbVaPVC0f6F5cBmStRN3Lny0HN1oFruB5lDmhVnbCC7abEHIXH2FgdrP/S1Ehs54orGYOG
5MuexFFMnEi+BbcpGTGt+ZyQD2cD8MTkInbj75gFLueAM3MJA5c29TtHhbYx9XyCZV7ti7fA59y1
J/4R+m0MssDj+TfNeBTt13lwPB7nfMPWvIK+fbiBDcm3L1YAWiZHZIfMufQJHfxw6993qFulINrH
+fHE6WWHsfTRO/qfYyXFMMxw29s34cpKs/Pgiuzz/wlUzN68UUZk74Yg5xaqfHMWdXF/OI/DxBkC
hw9w5Y8VJwTPsoUiHGa6SR0PgG2T/85NjeOK5Rb3ILkNcvF5+hZq+Cg6MqGsdG/r58wKfWjbo0Y7
TW83c5cv+2KluVxovDdvxBo297aV/Af/LxD33qzgS5PD/GSPUjjiZAkZhOM3ZLOzCorJsQ8f5aKb
Ztfq6ECmO1B+YyPDKE7Q65CfXaPYRez78vyz/mEasfyUXST84G/3m9N6vQccf0AsllnwxwUOIK2s
CinGkKTj3oGIe5DpHsuGvtkL2Fni92PyG9IWcGB6FXL57TgcVauRvTmd185DeSydH5zwBZ2T0oZm
uUQPgPIOsplEhmjpaN6JM+t3V5Vo2WJpqD5ZyO6JLud2Sylhzehs7Ug1MPdO0GksmsLVDhWBQfwP
rBUpt5bennsf/BwWUvSx8T1QZjpNcvMskRxMbNJnk+hdXxj/jsyFfQGbZIxbMo+01R8Kco0Vtfgh
OpZqgVb5wqMbYvrBOyllSxyJeJ0V7NvZirnhXXJO28JF+mTYoSD9QHIT7BGOwoq8771yD9jCEIYT
`protect end_protected
