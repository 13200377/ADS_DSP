-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
iXt7/J05ziSPPbcqVU2rtPzfmo8G6G4gPWdfRsyEho98EENP9RfzQo4fwF6hz+LdCY3h1GXeMjPS
6mMgC9JU31A3RYWFPRJ5lOpJfOWl336K6Y03SawfmR7hwpoIP4rZ45UOHgwPVUeeOWxMS/0sXZx8
G4iWnla6v+X/IrMaj5ryroPKmOEU7OTpx4nWGxaJWd5sxR9NU09ZHHK2nVavLQZgA/hoQUZw6Q4o
cx0YJ3zgVm8JlvQQLeKmwUqtqPzDfWYxXa0NanBW/6inDhB9NyVQryMcTvAK3AD5CaReIyknMFKR
u7rheoDkckCwMunjMG9YsJXan8o8ekZdnVL4gg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11888)
`protect data_block
PF4up/9vgT9RbyNQ40jQUsi29c//FCcI4fPtjbJ/Ui4ODrSV2Uu5ykRVhciNl8y034tazDbscNUR
QkZFeRYDePNOle5GNOpFC1t/gD5fLY/VBI8KLZVdSLChr2DFr8hDgNN5Ez9a0bELUPZ/NiZ9MFCI
bFp8AVotOCmoKQ4woV4htXM+EscJtN4IVmvc5xf7m+7G4Y2dDiXlJsPACrwCFNu2SVb5D6WgqCVi
FZLejuK+Z1iYtc4ywzZYsDKjEefaH9V5ZR6CIiWEiU+ccnc/I6lnB2XI701NlzFGi5ZBD2Th505Q
9BfLbhSz6dzq/qUWrDh4GNVup0ttnL4ooT7VtDbImYk8v7N6xIqRQEipPPYJlYEsfZRMtteFOmdi
XAp08Zo/jcNQ9Yp3vFReMsP9aDqrPK8oMw6R/1LyoMErmrWNwTJJJJzN/knuz5duNv235v2G7xjy
HBZ5pNMdEX3wsYnWRjoasQEWhOCecZCgB8Yhg/24//3eKpLK9pCQNDuzv4MM4tuWF081u42Eh3jB
nLgoApVONiF//e54OMOtSXDJfW9b8UIFI94zsR6lcsrgfyQcnLQ8TOj1bD5r8h//RXu3WjauCLE6
omNi6wTWaF+V/WqCAniVHcx+NUOUp7WGtPudsQdX9rNjJu/CQkwENhPRVBIli3y+y6yREcjEDlf8
hrVx1YighyJQYo1g4NWF9fzgcpLaFG975C6GTD7CbpMSh8MN9z8w+XJBh5bZmEVIGNddnHMvPww/
zNJFj+cAB5qmROs0a1RguUVVIMMoxEhozrvX8jOopDAG/psrIOiUzBgE2jqyaqW3bwzjSbz9ISNc
39VU6eBvrPdWE0QEghhGYGmR3ThDawVqxMFZOn3KhCn5RDVdV33XMdj7ESyhTvUUCUIwZ3CA2+mD
3aGhn178WhEgwMUCUIRiXK6tfhOEQO8xMJUMw/NMyDAFKmxTQcDUQQZSpkCPaP2LXhm/Z3OD5liS
MVRyOfvSx7/uWFIRipeWun/Yr38Pc4HJ9jfvNYKTRVd4fjosHML10AbxNwXsLUl8E75BhBl7xc4Y
ykSsStXQ3G8PIuk5ww2FF2Ka31nVdS9quNFdXEqqkJUUT2iO4a5pjk2FvYARIfUnVqMcJylKeKEB
/UdnM0sPvkXbe866CeHXnEbDQoEMhOUEDcxYsTjN5FrjYzFPz6Ciu/DF9tWvLf9PZjE3tKMWRqRr
U7ArApCx3welKfkkMBJ0vdv4fHzrjJZXjUg7M+i9dtjMkTTNdyMcGhN7DdeKfk4cdW8YB4RagwrE
bdmrRHNYArIJOUfCX4oADyBcj6qUqthVIr/EFO9H4bICivmoeHJzrzQ1ecND6g6maQJd7ya+Lpq/
L2tsR//TQdmnA8wUvWsmLzmYCaLysmq02a3CU56hiuK3vKuKkV8hbWUWGvAL2CPDWe/dgVsq1u4d
iMvWKgI3TPxW8M5ImAeQyWz/JXkWDxodhJhkecs42Pl+Q46Q8tAnhDelSsY75Cn/NP6i//s6QYqY
1DgMcJQMdbmEUuusOe6rxDnJfoxeJLFEGHYtYYsTLs77u8WcrXZNb5ZYpFkAwtUayQiOVQvIBr6u
wY9t5xqPIn8Bqt5L3JcCz3l+Iw2mvNjOA05sGB5AJXSWXJNDK3z2vBUmIxZUg12EMwyvrKEctobw
Jwn0qyB43n9fcW13HctarNkSIpTk7wQZYNMAA/g4m7wTHWZ1jNFKP5GShVTbTQgBlGI0dpiAdc4m
919tfapASk0Y4Xh4FCPh+Cr7UcWFXcG/Frx/eZKyi7xM1MEXb8JsX6Xgttes13reNLPrscYiY/ky
K9VQyVXyZr9z6uxN44Cg/O0pJn2SCOconpe9lbcBfGDaF7GauK7shSi7m/LiikzqgccDtM87fMye
gM1wubVqCROKYQmxTFmPZDoPy54xCx7gr9uJcLzLoR2NX6TVDAl7Tbn1xV6kT58cJrW/sMovy4Y3
1aM2KkUt6nbdBuar1tEFCJVImtSt8ESTVZwJDMq+8X5D5SZaXy3U6avuXKxU5ZuT0GI8lHZYwI3f
vVbb9SXkOk4/yt2/D0MN1J5/ADcWy5L7Zy6oIC3jgc6aok59/NH4gScy9mvgsaXIaRYGm1F9yiDf
WDlV8mfuyarnzCl9BV8rV1A+qbNvL9biF6N2MAxqIQmm1M/J4vKtX3SXr9jhd7uTNbpBty8GtqbA
cD0ETQ6+RCBgo4/T890Zxl/RcGVn1TKUOWn9aJZTHErcWsGLBqr6H7/VmEhxZslW7Kb3/i12fj5K
YlWsTy2w0995WdV+14rkk5j0480xDdg9hG9T+GU9B3wZMTYTVZjKNJ1rrE0I2jlA8ayYog3PYOFc
Pe8SbL38z+KFNlkfAl1gbexZn1YFniNSdnnTHintyXCNwHVcTBd5vpP4V26eYaEw+gfotFrZrhvC
tVAnIXby07j8lSOdd2HdhOHBqKhyb9UMDt5K8ALNWzYmBECKiJsZl7ElqHWwv4zG6tiB6Eb6/APm
/SY3CGkdwm7AlUxOyOOXBErADBs7HxhgHJt0adrKphbr9Fc3lNBUiBrRQZKb+uCPTqPHUzwfnjgL
85OfTd525YNtD6iJjW8mdNqp6F0AuYoGIID4v8q7hhFw1YhFKpzemvV6UepuXUvPA9Y3VOBIVLn0
VQe1mw+hYsFvN7BylLl0JysUU24nz1OnTupvymQoE4RY2rOJHn58HJIjlvG9LA32YiMnSbVYFkLP
SZpB/wxoopjI4sFCoxE/rovM7gycxvu8vXiwu9kgCIxrUxi9XeGfSLabqDtDywp/p0ZFYY3dqmRG
G82Gc32EiwEt/eHiCErfjMnh9dwlHWjgJ+M0g/gKt7v+L8A+cgBVKiYld2gA6/WEDgoK5o1gjFdS
dGnRSCAi5TXTcMY2mC6HXQiWieGBETCLZUeHRyngiM9pjUC3JgKbQUzx6Es080/aTWmLSXnph+FJ
W1F3F2Ubh76mshtdRTM8SYg1UT9FfC5vV6bsJegSsIs9jCol6JYVQcKXCqYBzxAjjxyc9cIjU/Im
mNA9UBvU7S3+cU/FIjO33t2isyofxUB/dcFKld9iZoSfjobP3tBLVGZesayc6OW1bq+ciMdmjm0w
r8bffQJgFQ4r7pWyI/KKqbuJZxefj14NurfPR69bllKJPfdef9yLXzo0bUAQXi4PpEVwXVZsU3Wz
96D3STu5O6NzfFsyv4Uxr8mcS6pQ663GXNf/O2tWUGqr/WOinL/nTxno0tV3ge0YhB9TW3sZIZq2
d2pwl0fzPFpHDmBO7ZioYNS4LkfYHeKtT/LJGCq4+5G8DIl3CVLBQkvG1Ybh8HaPQazbNm8aDyue
N69V4sEr3G7HFYhys/7jatkCByQ6avhtvrlJUMhzskDXsl0gZraHhIoKpgf0mClLP1spOm/ic10K
IyvrtymGvUwwIYwucDRmE1UaXvK0fUZ0qeBTSKrc3V6BZhKlO2CVFNEgXDO3JAoxAM5xC47XFlqN
gjW+A4SQwhUU+R13OqUbssL2HVhZKwwXqQ7Vl1Sz3ZADZuuVsvthNeNOI3xqh1NvL4N15dJ7JEmy
2aCNYRVfLTFfUjXtkEsVP7jWKoQzx/+Z7n3tY+VXwacRDOjr11uGHB+0LRUXdJ6EZxAIYotL/jGh
M5G8YRYfkPr/fHIo8SyCRsRoXRJwvryvdxCWndg87A0ge5VrMcF7lQP2ICkb8juvkx2o4Kn09Etu
Hf8h6FXu2PqWa3JhIj9WA0Ei2dP1RzTxR4RHYCOUb7q4VpOG5afLZodh3n5eG07iirD58puKjwjr
m3i2M7AA+b66umGmMWFrg4Cn6TyEvqugZAR2UQHaWMnl5Do9oUii7wk9gTItHHg7hcm9QGFSyeqf
PNhq+iWBHmJWXrjlsG30ZNxWtCh8PBa7zPRNS9l0airfLznfsw51pficqU1aIOEX/ocOlcGbO8hw
xQu5d5dvfdkLpTYxfIrrQPADJ5e5dFCTIAJIGSEWoRI9IRQ8bo3FIu1cUG4Lh8oTBwm0b7L73hqk
ROQEZcNrekssNn0NjAMZHlYSYkaYr00CvJasR/G5TR9ha7+IC18bF5fq2MFHJLfSK3K0p5wZTEp8
vTz3xH+FSojmJsQtKV1gL7refRl+B5UDgktGMV17efWMG0B3TAAd+2eiA3qk5dgs2foQPGVRplBO
43cmTtyBjiq936qUPaDG3fHF+HXwCvbkSxS91wTYZJfMWz4KMaxikmwRJb85m+d2BERc+DHJ2Hz1
RZbQsnWvytARNTx1kp8IY50uoukRaGAvBKaM/OArHhqgeRPkV7Zh1qo6vUV6eePL/btRrCn0tGaY
X+k7TVNUyGcnny0IwfBKF3PI/Ote3K8DJtdk1C4lmcW3EpnzicOv7g9443vdghUoR+Q/28iiGs/f
4SUihkLSKjX/spXjYSJnvyq3qTH3ZCUjMyK9Fn7t76YCcsghWRwJloKH97auNx0TcVeTGajfSJLL
dhkj+cRjw4U1ufQgjpPWwbx0zeRUO9LnZaUsP6ppA2ToQlNQpeEKbIt5OqxgHDZAlOPeJtjLthQP
rkgRrHQ3VTST3AYho7+WkRbJFlmlI0Apmte9wpSqzcGIKg8ibqaIy0AIO0R6QbjfG3P1FyIVYzqA
OS5Tv4ghIckkI5zdM70Lf0ZHRHtglapkVedXEVfmjobk8ObpMlVgcy4uEdJ9UZQSp+CBKemZFErj
fHO8DPk0ulyH9AZnXNrp0IaCsSyGB5iT4jP9/00pya1Mqyd3l2R0kBGuECvVWyGOY8ORef32GCMW
bFcXQrljFgpc8P0gbTOMiQb/D+qsgsFVGLju7ZUb/iDxRsk2qCtvFnhK5klQbUCKsV7ypM0niWLR
v4dti5IUyIIyRY2qwC+RJXMfULKZoI/BseTWMvc4uSMq6GuPdI4+2gS404FIRX06nvWMU8QS7x+L
GsVByKm4ac5TgDX+Mu7IRQMAjqiOP3Dynq6HTfTlQANSe5HdXJTngp0fZg/Ym7d12emZuWwCRz+g
8uXoV5FYKd568SM/9b9VgE47ZPQOdGsJkQA3lQ1UhbgxOc3fT0S0PIC9ew5e+rVdK2DAfY4gebnZ
45LsOjWSDERfGrnEVZEIRBOJEkj11OprtWL0c5gBPj7ceBtzrIb2x4E3mfndagHNydN0vVF9E7G2
hgfNoDbWOq6fVIHlqxW0JHCWMaQPsTO4jYKutWQ1Y+z06KKfrelgBTfwIT9k7pVFG8SsPSFcnIb+
+2mjAFxvKOJo26VYprHVXOT7ogXK7UDQAfyj3fnP2Z8A6DR/LtO3c4SemEqfK10ekinlEc2rWS93
HE15r85giOEF5buxkm3RrC+IjvDhpj4hAGevhr6VpT0RvFf5oins7L8llTD4SJXKHhFVtxcu4RS6
kbwNuPvgM8eR/N+10wdIZVJ4esPuqbPwKkXbIOJH/S3eAZGXLp9Mal+ZfKIgtXVa0VWaAllaI7BD
9c/8Z+oKgXxE+vhgs1vvpK2CF8YwWNzpDxonrqGQJQmhVabyBQLcxyQDrrXXhPkC52h45Ps14SDm
qmOAh2wgATaBIUss2IP7TNxt4QSCdwqVzdlBMXc24dRjE4rAQsBfYifpFPG1usrSNacBGm14ysKj
lxcWNLiY8UbpatFSUlnBN2PJhTAOeHICaUeS880XQUoGIhgDP8GiHzBB6An96dTK7AnWRrRV0zxr
ki6LhRmh+iZ7EPx5UVrxrZEXM0eLXrZ4j4rfLz1Zo5LgCSSn5MR294mPBvWNJvxoLzzeIeQVnSLY
u35zxEykhOgs3+F5uotIMlQVY6hjAZfnNu3UH9KQjp5+Lth4TziTSfF96MxvFAPIyT3qVhOdmSy6
Sv1fXeaRkwgGCRres6S7AX0yIwIv0OvxWvQNxhryexv/W5BGeZNA9z8qwToaxgN6XiLMmFhFNXe6
d8xidKbTIYvnmYyx7gBDDSXmmwTZ7mRqJM6bSzWu/56m1u2OmYB3vaL0Rrmch17AwzXx9ox90CSM
WRzSRvEk6gqyjDY5kiPJRc5ojBgcbZKzV4w1yqF2cAcGRoSo1dJiRYdEygJ0XmSJ/NW29PWzS63x
5zvvBPPfuAOdGNVZdp0oblIW2SyTmYcCxW01WQmbHq8VA+u81TrSRa+ajIZFyoAGoXY82eX/Wwam
F7lRC6Ks0hYssDS/p0wZhtzVp/pdeuX4QliJUMP8LqlPKiKFwVNEKcucQKbPdhob3zj5My7d3VrB
bCKl+IUOL3aVs0iIbgtMFA0aDTVpOwVmteRvHtMizTzZSWPQe0hnihRcGPRfiCzz6LaamshcnlnJ
Or1t6XZbCAXF+52FlJg82ybmc9tP6BkZBBt78usgcP/I9lxtnHfQ/26gjIdT+EypXIx0P87iN+7B
a6jJbaWTTAoDvI329jHFKjqArU1mvRZX901UIWzEH+8LbRWD/dlT0W2wzqDNIin7AfBBC8Mz/NtY
Gy82uJ9gEigdl18vGoA5eXE9jUnZFCMz6NlNZsjDtZlgf0qToj4YdAB0Q5v7rTsdogHPg/a2G+O4
BX4T4aXIP0cieIivtRQ62fsa5bdbZbHPXBvKllTkZHikzgjWpYvB3P/PqAg1OvUd3U0X1exVj5Z/
W9ZOkktMnKhs1hXgX6/Ev5Hq76ldSrXn3CWiWGWURMECLQ7/2gGQiGeiqjLBzq3bibQslAvPwElk
3d82Amiz5C/IWyqZXS09lMZx43lP1BZ6W3XBWuv00R0psBkZRAA01nXESq+yPiT967ZvrqPjzQxs
WMeFg8ZzUqRQ9D1PsepdFwkdqGjGUExhuvbO37KjsFW+fiPEP+GFkA8ouN4k/ZtjOL1ufk/iNj21
ocnFwOd5X02URHB30SO5Ag6zzvqT8JKFejSaxAHXTy6uEWlbgcCXsil7DPEtzUXbZCa3wKduJdZy
GsnjsmgxXndICq7imEB4BUkVwdMs6zWdkXeBD57/hXAsCiv6QpfrUy11rmMduhVaJLq7Lgbt2hUG
Crp/L5pjUlnDdf7CHuit9U6tWbkUNB1lyE6xqM0PSC7LvbF8t2KhyhBlo43xPUMo3tP5+CDDMaV4
qtgLPf8NGKL7YbJCUG4V5Kjv9Cmj2smZg7G0XsARDTk3jl0m88SJRv3p74MNxvILwJpDxo8+7L6f
OSn2T7aU0oQxCs6EhFACWfBce7+dW04WQB7q25IE7upRr84qsOq81iJA5/HZkk/iytSq4VwfC+UV
UH1Yb5qKk0KExeK5ZZQIC1vFYxWyB1h1TPZIMk0Z61i7LbCR+rGXaib6dtpf/Dqn9aLb/GQOi7ly
43esXAfyy1j5m59Pb1FN2aGeV2Gwzs7tTHzbbXYTJEnk/PoVfJVO5691ssUGvqyKFGYUC2+cIdCf
rFT47SCRcR01THna7ajDP5BZlaDtc+ujw4ItaVBSXIi86o9oSjfT5NrdUvXcMvNzcpAHTINW7MHp
gDpGbDGv6Z8Nu/o8bk8YfJJ7gWFEdVRBxVnAliDIrRIAfAYhOtcKZiphbVkUPVUqV1CF1XpVfy5F
TwXOFopGgjifudDTOl6v5W+iqMkiSfPJ8Mha1HM081hPyv2D4bnmQ7VDIIEavay/R+JK6HDAzXi6
eaeKSRyIvybYmMpxufdJz2x3FStIbTNhsuPoH41wWqgiGuCv05eI+sF41Hu2I8fPLx49qmD8WEM7
Is0QT+Amjd5M/sFgG4Bgc4RxgqgvX5gkowYv5GIpMCqI2Qq0nOgQ1tIEntHuxvopAp27gRGuB9Et
eZ8Lg6vW5tekSw5PJGWkInCyCjFTkheXeV4aeGY9SCODGHc05BkLEZYmjgUlffB+X2gpkt/e+CMj
ane/BqijGRWulYpmQeIOuLYd7wIWGdKmA5+F+q5wcHKolO4TesaeyzlvQT6lquKG33YLqltnza4e
0Es0q6oXfl5cLtDr3O+AxMQndbfaLXrFxrUgBb1oP0Vx6IqDHyQcplZC2ZTGBSZBhmoH7DIhsqM8
gP2QCMEbYMAQWqa9Ccn3jC3HVGamGDbqukcVognSNE93OnTpH9f5i3QFty7GnHbPGTNrSKbcUGfq
X2qsxtiCsAxhm4ruCR46FnWnn+XDOQN113bdN6mS/sgFr+jy9Zcn0rP54Tt4AdXe6OB4emv8pj6b
Xd2RTcw38PIiE4YVqpYMAhHKteh84H8qsGt1pNobWXkFKLN2tHOulctRynX2NAwFPsO/sbP5/UXN
7TdNRnrRd7uRXMBy5Db17TVxR/gaoe92lrgRmxMmR9zVzH2VPkD3q4khDY+FykhlvoLXgwJ2aRzX
qqCpOjJU2yT1D9hgjhKEFbxPUnJ9Kx5LOv3X9pc7dRGoTmVVUnG2pkcUZeFfcH0e0LU6EYsYWO9X
Ymp+9xi+bQ+fGX12pjCBSFXS6TffbkXWJuWgWRWVdSjhKO4jN2fswko4KRa9WeDDaxBU+kDtpqLV
CAo0f96896XMZJ35VsJ3Q3IozJQM3FW7Erf6r34Dypo9X7R1q+haG1S84OAqAjwcIyDZSlnktmtB
QDA5J/BnjEa3EkUu57VsWGFedEIAmxN6s5VSjq9oRfxwTe78sWS8L/QMb+7AByu1L5KkT/qqE/BN
4xqAfnC3rkEgn6nPJkKmOgW0YqvWPVJ34tpNM0Cslfb1ZkWZrRW6K/c1RlppzPpjGUem6GbSiavf
vzL5vXw5muMw1ZmScRXXoYp63X1rWVZQZFdKQAF7wihuzl0/cF2/plLU7xQJSyQQE64VqXyhE5fM
TgPuXDTgssidqjreZRlmy1tlG7mJLW7B3GjCKb9gPGNh9HDsbxBqrHT9maXrb2ColnddNvG0UQTv
5Lt2pzEBFT69c/LErIsFy2dnyg6ZWxL5+UVTqdW7CPmnqqZ8dwZfl1LlDHyOwGKBn0qZowXd6vs9
pIMJxutUxKK5V0/hApqz+ZF7slDSgIrUGYjHye9EppCKYue9zKzlcoczm326GI2UWElErsG1UZM5
ihEAIa55ExvkvZvHe/rACPU9/aPetds8s3c4G72q5pgEVcP9wixrbfgYdec52yAM0a+HuUQ1/IQj
JFzG1lpdL8omT/Q5UFlAMDzvC1sJpDZD9jHXAJ/OxNuFGLbPgKM/gD/KwlNQpEqfk62yoaTFg99u
UYA3pI8ZSoxNiJtSVEqGtCzd0Hp6JohmSqjxFiwUEmtPItioAHNytnx/RayKPQTFNf9iLMW0DFRd
PR4+zmaMDX3RrjWA98FfLLKzYnFDFe9oBcyeVE/ySR5820s1kGf2OIWZvymP0xQdfH+ZsSs68Tu2
Nh7GhCgLuHzJJ+RLNJhXQnquFTKqXIZuEI4krgXghiO3PVpx0j2BZxnW8Z++fBUc2zGGnw7DkUfh
92T5ze2zkFW0PzUQXvplP5l4ftXqiTjlBSjg49m2mXqXgRnzPHmQZ8CLE16OkHn+YNPASlhJnJg/
jTmmieYQBmhFY8nA0+vIctMwARmvUXrtZcBbxh38Zgj64pF32l5LQTyf4CLtU606UbMNM73Jij5N
VgGfOp9OlzsfrS2CuRcFNWobtM4WRdQKZjV6yBdfdx+B0n1KKw1BVlm+mCwCgkmozBMCxdHfjwVt
pks0M4KMmqR5NZlo05Q1LS6Ry6DNBTBAEJJ+Ij9QSgFtaxoQZWXOf3B/TV1+SmJimcKIsQXQ5x7T
5W0TFwhSMp7cdRY1ZhHzeYInKWGfVOX7bfM+yoehF7k/F1jWEXYc/NdcpybbZzyjoHyjFjqrb1nl
6PwEBIa6ZuXPA58p+uD2OH1AarpwHb6a9rtV/ZRq4SN1DFazRUW930TH9B5St9jAU8t/sQ4/KgPu
Xjkj4vr5qwqk3oKlA9cwreh8A2T740TxFspocLRiMT8Il7Bs3Q2wP+4KnGQd2rxs43f9L+58/Lu7
rvHiNJEhLa8MKAI3ZEraOlPmjINgwQ2KpkbNlbx8yk3Hm6oifWoJDWsFAFXw4/qAxlAWUommKtth
CoHYB887T6AhWvWtQLMXW2O/g96Jq8p7Lw+fP8kdBGcX1XQoizQLRp7+4sAkeuJ7vNvTYkBwaRKI
9Ome0zd05bubEmKOhluKtXmS1fEdlUTMblAvenMSs3XOMXy6/upvdxFn/i8KKF/NAciu5k1LqIGn
v2o8W3QnSMl9Amu19PfvKPytObayNlQ6/YgO414oYt3XkImzf554rOIKO9Tl/Y+unlHmDQ0ri4GJ
rQPxNQATAGTFHc1wtuBQha15I7yeVuj8OdNv5yhX5VwsGa2mZ35oxXHJpzyiAn3WagHMHliS72pD
lA9NPmyGJ91k0r+qEuRfj9AGfTlgQyJJVNqu10LnGH0qsqdGZ5Hrb13xcGgcNprZlSG08LyQX/cI
nS1EjTI5ZS13t+R6BpaQzmPCEQBddhjLDrnuNAp2vogY/BU4155DPzewLvzQwlvCX+gSRicinKdq
VWV0lnX0EzvnUuJExKeHFKdQ+D71p8TDVMaCiIp5Cu6XynZChuDBJJNPIBEHqHNM2VAciAPxpcTI
3zFfrdtTBZRHbvuSRIWqpSLg4O+Pto7dYZHVhf2Pc6khqZgfU0Vrm3sKlDxAn/J0wmf6jKggwVF8
TIqDcIMyPyWHf7iTxxS+jYOXCjLhbbIBABNUvWZ5M0zYhRBtF4wJ/wPFgUzm2Uy5yAIf3RQ9uiqD
0qZkCaVEtW4IgQBgnXgi2ps+zZKohWD86Y44yDOac4hBroLuEaBa+0xjb120Ezbt621klJ43qvLi
G3deh/JCAVrxKtbaq67cr2Eqk9hHrDnyqk+Kgbv+ZwWqR7OdRApWsVDQ780Dbruc+HbDELMTxuR4
2A/iWYSKhqot19Ed7ZSVuicAmaC8NL9f3ILFue3ccWT7gWy5WKBGddqy7sQuuOVfD8EutfuyOs7Y
MonRGB6f3CFVIk2sRlRh2UP7bDVwMAL/MHf79WiJl5Mfx/8iVKMqAyX8qkb6DiFnTNlX3bTpxtdK
LzMIyHM99VFRYHTAMN5LFYMDH3AS67nTvo6kjR872Knwsl+M5WNLf2K7kcJpewUaUvG1ajXGUbkE
TvH4kEDO7VWnfxgFTd/yoWDPml8Ix8bSTkJR98xe/4mUvAHpMAHDf3HpHeVdS1gEoz7VM3KXTlzL
MN/lKNkNp/x+leb7atrD1noMpXXaW1T1b6dPozcENQwI7FQGBlZBcy8hE7JjkYpQmMar/0sft7fX
/9n/zDbn+bg/OBdNunQF6wvitcgPKzMUZFfBdkqM308QRet4mT9Atx1vcrJoZBoXcypGNOYS0+nY
XSTpyb1v3Y9RdyG5DHm/JpgBcguW1Y3HU6Fed9WgVAAoeGYOzYXGPeNE+WFf+qQ2aS7xjNd09RBW
56VfXfZjXstwa+8NyiVlsRcg28qPEUOpZMz7QfWroB4RGY1oWJd5nswZ1/z2sRjLwHKWnbgH2Jht
QgJxlQuQGgNkqRSZyv5Jmz06g9npeAnsTvKOCe3CDfTiA5fm0Ta1nvNbuSgTrRwjabBXmVPWIlxj
mzkys4gcOzNVcRDkn6/ptlveQs66CW5j0Bikl/Ek3OlQCPCSWXQYbA9DsaZWDapv+5qlA1iVUi50
JMn3kcnJpqvAEF9NUvpigYMnhRRl6j6lLNBfk5n8jBvJmzlO1h6Hoo3GnHJPq7q9mscR3Dh3SuHf
zTN5rsdxa44mC+gx+WKc7BGc+Gb8EY+HqhAszeio0nv72PH4nXHIQtZ/0EOlF1MHCH0Kgb1PVHrJ
hQBBZKE64V3ez1x1Z7saBErNB+8hMA3ZDI6MbquB2aT+cCtzi1SoHUmIEII6KEMn0Cz/6Exom1VC
2KmNr2we+ZSG/jQxxUCTN0ZGG5KDtyMicbaLQJ+simtjdHcioOSoa4pCwFsGifyU7j97BAAOS3Y9
30ETCVzn59ze3kG5yKHid4V87sDRL7b3LFmhRYY541hulFDucFiwTQ/7NHVuL5wTJBy5nOLLQVlS
A/UtnH+ZWIuN9xLTY66Ub83AbB59fHDiKnfoKc3iYAdqzWc+wq7/qfFr5b0is62kyMKHN2+hd+eZ
RDcp4eKM38eNuuUF+QUt+yk4eG8Xe+xxwmlZmD6u9ielpGg19zPEPqmYmgX4Z7BOynHflYfvHBW7
KrrBwxj7PO1U+R1q9InxIEpqCb3KMHIBsU/3aALlutS7dLMLurcn206gROIs1BH8krfNpf3P9ecn
4HhVBHkp4I/+plj9TF3cmXapHziwcnQ4dK6kecDJx3GVAptYwTO5l7JiKtIMPD04jqsi9EQW58yn
Bwk9//Chn+bN8u1KKGIEf3A6GDHFZGzWAS8+1Nv54zdXsrpuWjqVN4UuAfuC+wGFj5vTTYI/TsON
G9d/dxsje9c3dH+fsBvz5nRPvJL2cJbOyEUeppGaCssHnehpg0U+N5QkNIW9nQ0c90Xj9x07PJMc
NiK+AcqnbkGK66WgLxfnvH/jQThZpGcgD2rVje7MYX/0rAISySXih0MglkCR6l1MKjYneoY+1lts
JYzbwKQvrgmwfUV0SAEg5qLZU0ZjSGsNgVdnMXj1aTA9a3/XDp9BQ4ocOklOJPsHQY8lJOE1uD9S
9KOt9D389IywSG39wMVDDIu7cMLk0kHOdG1ex/+50OK5p3ZzH18TaBHJx8+6ulU6Rkz8ivG7agW5
JK50X8mR4nKUGyMUxDNI95yfXnm//wJF1iaG+c2jSyk6NsWY37PFPQuv2qbkEXtiuO3c2dP5XI5I
t+dDfUchp8mttomfwOh/d3jAKUS53v+dueu3esuxxOA9mCqqnb8OW4TJ8xf6KqR3/JfzRr9X7BHF
LtBpqPsh6lVfFD12yurqi4ayhz2e6cfuxjWqh26CIkg/XIG36GvNyj13kTtjrpiOh7Q8H3mOszTj
iiDCRDPrENq5elGbD6QXozxiVda5Xnbqe/P7ZFYa819dYjgIzMY/aoRWz7z2XmvT2kJHiZu5NbZK
qIfXdgheyx78wmwD95mdiS7Sk0MnPbUD4hSxXdxe3hE3YHUBowgfyItGDGIbjXkRfmVfIL3R0TEC
QE7bwtP1ZPNLHghy1EimDKLPEjOlyWmdSEn9OgPo2/7MFJlpzhnjnOc7GBAnKFTUx8ibKBk5rtha
wjM7b98E0msmu4VUuAIhBH56OFpRHqbKxMzOLaHcEKbZwta06OETuNXZaur/ai0aegw7p0KuThfw
8+qUSBsx0IlmT1LU0XJvqwqpUgNWfIKXVTL2v5Sk+AT3YFRhIs+prN3k3SO+yBPmB4Gmz9CtFn4K
py2Rb3nbUW/8rZV1m0aHEAmCSRtypRhTgXsTJ+41w1pzqXvIBN1ACxEkU9Ps6YFCAq0ylQUnmxI0
kHJ+heRxOgli7mz6QYSVgsAbtcICeJTRb4dyTTgggH/9Z3zKMAQG+9pPKCipponfXrg9xGC2mluX
1Mqt447ttBKeZeUNkc8/HNBB+CK3QPnze0kb+4oA/wP0hsffn+JpwC+6E7mEJof1czFtM4MnldPA
lsElgjlwa4m9iEjwoE6hNR9Db4FmvCRLP+s3hKGlkc/fGn655FbGJcvgVWnhqj9Bl98l9mDqGqA5
MZz0np4wIuGOACqfJZI8GQMQnEYkla9ZPu511ACm5VQ13kTUNmaGlvAO4iS0UTLIrmnn0uywlLmJ
9Vh4V2KEc3F27xc7saDw5YrlBFzPU0dnvJqBKUf2nFxwzsjXnRi2LrIXKiAbT2WrvHhTCWHse0qm
VinGSWf5A7rv+ylFtRZPTIV8P8ZWH3fmjZHfmrVw5etQSlsrRD4fZ1XE5dLnkqtCC3ys/cJHZl6X
IjxjP51ayP4qyVzg6sA1RvDnXZwZ1CmML0mXdgbqu/CYwM1ZGg5svWl64PJ0QjjrxHLP65ltvFRl
hrb9EftegUUorhzW5cAUf/qCE+Mefwmv0xs5byrt804G+bg7ADuUeK6YpwCbCN8cXMoBXQG3rHA1
qHbJP89ESItolzq3P44jxm+bQiMCGZ1dXocrMZI1cJ1RO21nvrUdM/mn7xtS0u+oamOUPZ8BHNnj
09WfXZ7BzmLTqjHtbVre9wvXiSpAUDrQP7B0tPQBkj+oYhKC5XW5fny6aZBJvRL3hTWDjqepdr+G
0090yb2jeYcFRbhJVw9L7GjPJeW5+xR739GmCuDLSWRdZBfkddyiFQwy1iUofMrkaSEVhm5Bbf0O
M2wjQ4Y1sbvPe8APUoR/FQRIzkW+MrXky/CMCBY1ZcYRaBai05Xu6JgzlNdJjHcWfya0CVTth/n5
Cr8d8G1N33Cb/EbKPVt9BvXkLr5JUq7PILDPkFXEPoBuHmi52VA4yBh8h3iev/h0lAg63mNBtIWW
k3ICY+FpSSg7q0ZSBxwMtw0N1Ud39MkvnZJOxQ9jWOGHpRTxhwMTMuc1wsev/ShCfFJ6scVTKlrV
m0AbF4iYmd0AG8wLIRLNQvdq/cQ3Mz8+HMJ41L5J7abA6vwqjuk4DmxnhNgeem4K27l8CwT3t8iQ
T54lERsmkHmBsfZBDbGsyrpokWwCOHEZlPc6C5qZqx2+6lAvlh/3AWmyHXnaoMAE2p6D7HbRe+qX
1NY+Jf0mfNSTIqhj9M5+ChF/z6ZnYE5rUygX2Mwsk2Xca79+OgthLTY1XQxlTKmUaf1XOqJuz/1T
ew8d1fVcwJN9KdsD5R6qE5nc/nrX/uZ+ryNS1I9LchVSpIR3fBY7dJhm1ekVmIjpVyLw7oP6K3Se
ikV3rfyWgtP1OW8oIqVDLztHCHitgtV1WTrcr786YRQ1WtjuyWHRtq/nA/4jIrE/egYnMAbJjoeq
bhgPxNDIVXwtIzzwfgJ4IUjZ0oRduL8Nb2HqDoDj/3gapkAam4V6HXS894nxBTTvlFBjz95KO8u0
QZ/KMBiEAfty0MItevfYO0ZqxkEDHlopy6Np2yMFQm81sNXV6bUn1ixvoEcYbPEL8Vkgk9WaoJWs
x5MncXdqJnXt4De6cJ2zm5x/ds5MeGAg908FXFjjiWFUv4OKOo+Vq/Xrs1O3GUNpQ+28LjnrnK0H
cj4vaq+PZMqjY4bqnJ26g+AhWH9Tz3izaLoVE/YpXU3MaHmq8zxUqnhcBRF2JHcBCsDj97bHsH0b
OHakAz2kTvrWio4Tb2co1aB5YoErM4ngjkQvrqix8YFxN1MGha1l8QR4bm2XLpaZ6MJyLGFTFkKM
pXZFTsFFCO4OHeo17T3D/BikT9IQLhKdmKBZ7B/PInCCLYR/cFCOj/rERUOIGMHL+8LF+Zm9vPaB
rsBwiNRqZokXUwRsAyQ7dr/A6uCbp38R490WAI+dW0FIWoMFJx4UWgEj8t8JQZgBDpXuXTuxnA/V
ZfSC8ZaUK8BiiuTb3AMXFAUgoAATcBjyLWcU+c9RjFaOXY1BWxOubugWbXQ4KzST/AfRSI6q+DHt
3sK8Wcs7/Euy7JrR4YtFooA25hcaa/f9WQVe/3G4/+5KuuvH1RBTnaA3Ycl2usrjbbt0BGD9D0IT
d5GsefQNxv4OO2XsE4/dfilRsiklbGYKd39qsjPkCs0AxuFas/fY5nsWgl7kSU1WIr3ebYMXUYrl
ct7zfKG7pcERRZ8kzKaWTlX3NQi/rEcFZHpLRMwQ39I1szQjx3nwuuMAvPx6EcB0IxLLIE/xULwN
+m0WAIVbP067Xn3wbPnAuUUz33YOa+ccDZpuBjWtorsbTFdnO51ntm4w5ubR2tp548hIjZAhjmwa
bUBg6NrqEkRSonEd9UMdWfKIYlI2YkuTadRzMu25C7ph1/m1lSmMa/DyJAOYUIM2wvmOgaGUd9lw
cRcoV31XJgpYbCrQIUXRg6qhtGq5dR7xtpDM6B2N8oLsewd0rDpOaX2l0zD/ZA79FRaTAgUnZwUO
eSERVLF9W7Rtf7+uYhVhsWlg23kp3qoa7J7FGktuWiM=
`protect end_protected
