-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
lG0QnIpiRqkauJoh+egi4HrsFjZpVWJ34l/TFXbyMbiAu47Wsw9T9KVGVFE6HykOVqXGzQ8lQgGG
c25gxQVfqL53U7WMk6wb3jNg80MArrubmafNNYWOpCLDyZ/t4KEB51Jb7X6+D4P/QQqYLlh/2kkf
oKBUgGVIZmb4jrLfRViMoE1z3ymYTdqO1eIG76aAiLvhYsvSPoFCzV5C0PR4HUwQvxDDuF0e+e5O
m5U2BMgPJjqkpNI5f7AoCAG4OuCC+GawB8alePOXCE2KaSsEeq1B3EYTkfzB9nvnXsv2/EbEHRlM
bl/fky1Q8nrNOysBV92iiWT+YetO+FwgBFaTXQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7936)
`protect data_block
QOHgejhyUO/wbi5myaLQr8hP4RzltJyhPtLE+r8r6p9EVT3+3N/A6+9mgKa8h1q1TzrCRbzC5ouf
UChhOJ1gPTTryGhmf57y3T81j1N0tLIRSmTnrXjJQVW5WikAcsg/B7P21p5jso0VZT95d7+m+nBP
flxO4a/va2RZncfjrHWFd2wRhGLf0qOqd6rIYAcueOIVCE0wPwoZuVUQYtYt4ZEkvw1qTW+UWqc9
LRwGjZC/qk83eus/Q25iSemleZCiErsb6dA+wcy4Hx+CxOJFiOuZYOSVJPTxeXMrZ4HXEhnIhUZ9
2au3P051flfG1zy3HzBIW1NfHstst0CtqTBtapRgvhn5aLbZSVrd133Ao3oNVSOQHnXiuRsqalj9
PXfziLLdqwiCQe4OdYZNUSKI8i8ezS5Ru47WzsavAoVi4zXiQM/O7/DI6NG9CGei66rwWS77OgTk
5z5BOm1Bpt6szBdhp5Pkde9QR1sgEI6tuX7YSCA4LRiLeP8t9CJy3+CQvkFD1APKYoxOMcm+CYLy
ISJrcKG2C2eRc5aEZ9PRpLF9Of/hiW2Q6kfymneRUP0qsr5nAYOa944IPgtg3VmE6DUVacRBtTM1
C1J/3Qc1iyfez1nakCG///gnXmhluCojw2fycNmvR/kBkSuay7WOf4teYDdSn/nlP4RnmSwdC9LI
ShQBv0ymBDHcLfNpivSpKNgeFmjkmZN12iilqZoGRMz1LrZNYstJBssvysPQlCE/KVkNnmR6hTfk
O4hTMBa/SQQxtEPoe36h/bNC+/PTgFfdimJwED7RFhNm8Z2yVIIFUIpAbDGVdW6p2UkpE9go13md
Bob75Wtuqxkf5l0t0tFOHgkgRK/J81dlfaYU2k81Ky81pp9UQePbitAoA9edsKgJbUJy1Wpm6wgz
YeGHdoXNlqZWJTOXrKeMYhZ2fkrcuyg6pk6WFHKkUpTSBfubXyds7cJlAA7oLeAxqg1GkbXbVfm7
LB6UpwDLwR31WnZpU0wakOr6gaVufElJyLTWMukmt4EaA4uxf3zHB6lDT9TZ7gcy5Z9YTPYf5+T9
09eTrTB1x3N7P6Otpb1vABxGmZJ7/j2tqNnyYONwRKUZWvkcGwoRanIkdt7xEmctk7hD06s8gCJr
5JnVqUr21PFfYw8vJVbFobUheGpe8ctX0EGAjmSLsDFEDubJ3RzYI5z8sxhHBiSz44UxDpPCKnpN
xLDJTwxP1bMalwOcstlzG87l2pnQIxiFIirfK5booX/S4MOkjCrJY0sbgpvHiVCOq96sxAseo5bm
M8YXPAdB2WIzMrwtcQWG6E4RUOVTivbRadKJSn4UwUTNvPXmSHQI3LzxtxLe2uZuygMprY6Anz45
iP+lTJvfu0UBZZcGG2+E2+2TX5Mij7sw0KjByWlNV5p3EoGaz/3FVe/KlJzI21xevGRyOTxopm94
XzwdCvwNOLayDF+1xSCo31GbgRNTfEdFBbZi2a4n8VcX7YUZlHeROSCxEPRF6o30rXLO+te4u+G8
iIwP/RaGwZZYgJzBTvH1VYP0OTo48ba8D73yundA5IrgL1eSLwXKGvJaCrdyqkDtPLUof7sys9l/
5DIY3xygSjkuw53bZ10EuSqlr+1nrg7/x2RimHaq/1Drsm8t/9XWORrXrSAayBNGJkDweztUT4bP
1n28AQDNJ2u7X8U0iAxWwq+kJy6y5yWi70z/Y9W0eVWD/9ZfPDT79dFRsibKAcAae+AuP3Lnwu8T
WvGWh8QR5j/wQronLEZAJO2nSphUHJgCKQdmRGSrC2r71goNCwmSj6vOjyyXXwgmpRGhZ28e69Q0
2qpqwSzkWSiXd+07z9BKV/2QWYNU5c8JMJnkM6O/9kBzaRsrEIF5FPD98FL0HYQJvx1Z5TH6sDxO
D9UX9flLXc2XR2ef/DdTUZm2D0cRLfr8ClmSxQ5hV4f3L8yvY8+F1E3to4GF4zFt//xe7sBvQNck
wBwhC0V5VSPLvO7v62MIlvOsF6SW2sIAExZhp1UyURPVK62usD+EAYzfIxWwZMFTQa4/yZcMAsyL
v96NBCp2umIbsy8Usc9JKdKPr2expzsIQUnGxplDpPNueT4/6LqAM0Ca2arga2ZJLspzxMrbV3NI
rgD0cYjSe+5JYAzwQtZTQePkZJ9M4P6e9nV55oyl2Q9wCbtlbx4eGJc5AO6WqG2M6t8aIG3FJ/7r
33zXLXrE5gg0Cm+P/3+edGNichJ0xr3HnhMQcwv8VhiEBxad1/0kwMj7pY/YKMoKd4M8jwLtIh32
EGjP9PQzJkUyxgL7e7OCkT6LIcAhUUfZoMXQBIn9IfemEKduB8AS9M3+gKxhl9qFKt+O7foDsNKD
s3J9YukzuBzyxAghxMxK7d/bD4rSy55asCrqJ0TdMUPRp3DFZmH2O9WZ9GVoy3toVc9XSzva2a1S
Q+LBwOjjZcDWGNRffR9Jn2vSVkRcSnJV1nRhePDJ+JMo2FN8wk3woGPN5OMtzU8cPJixTY0PN7ur
dHJYWgxOAUTR6PmVqowyj5ACa3SADWezSrnX2berjqlxNy81ofvJ9dtBdKFxFrQb2Nhtb4QyC9TH
opxOHszV7VxoJKUlJ2YfKiymZoRfgzyEmJW9ahlE0Cs5X2fcYclQXLi8o1qh8LY3a3GFYy4W1Qiv
Mg0A7kyVCPGGNYsFCXsXmrAdpWxecastseZEEnocWcP9e3hnKXE+j7Kx/u1WzC6VdhZLHv8REItH
3w6c3QB3JauAhQSpFCPZ8BsevBIoN7mezT2RRjGMQFSRrvd3qtzxeAvdTkyfjgdkV3Yoi1UW6d57
2y6R8g7iGLljJSNBjXQTlTxSKDZGJF1cL6x69w8uRiem1cDsiMi/xhuHoRKT+5wtEq7XqfQiRb8u
dSef2LT4kyz/3Zk3RIskYIoFXt+xarNPgtfUVQTjtkH+4ScZgWZG1KpAw6BWkKiqFB1RVwLOYjQ1
wrouxg+Hgx7ua6F6+0VOK/Wo8sAHmSIuBv60dqei6kcw4jsWhsoEjl3pllhLB+dh0Xu5nFSx1va6
jPZoKP4WVXX4T/vJfVSfBAp4FUf0JmGEvHMI/hluuY/vEDT7aONAjY1VHYEPQILKZFsumKq1Dzed
1uTabe7/t5+Mw7WylRIuPSFs+OrzHi+qmrT31VOecVYBkuv7IYSbXZ8kozqdnJfBIDh5aczlcFgk
WqnK6dnZ7euetfFM8shWxRT2btIshKTKXVCaoNEcbMqtzn2xgy/SbXH884x2fJSdDVHYd49hdSB2
HDrV02Yljag1nDCg+8Bjob38dKj5HqQK+Jhju6kWfW7go79rTG/fn6zzZPUwFKdX7syTmHYpTBYE
sAqYZR/2rMqCMnf78kTVxiwIVWu36bmnh9ku40z+6LIiC1GZxs8JocsOX0L55Y3MEPgjF6xyehXw
2nQ6MXEnKFlrcAyLWGR3SpG8YpLk0+FD2MSbc5y6LW399zKRBdfl+Dbx1VF1mpkDt+Q6QyrqRpsC
Hw3LgLx6kbLDIBzObPtBf/Dj5CBupd3dadMYaytRohfhQhnOxBcab1DcTIHF8WxzsM2Gw8ZTniCB
O3kPGeB4zhqIN/DcZSG+dJSqmyRvbWjVGlmyw6yhM0nEcYx6xa9ZdDqvm9G+NJYZuML4WjBBfwPs
kj78h6QXP/SlYXbNeqao/w/J2yDEzgd8uNdUq2AGxJDROXcAoDvxkpWNGdYxny/RU7/4SsPvJqyd
LPQArmUiZM8g3wIoGgoLhcQji1/blp6eAaEWeA63WAJ5aAQ9pPihYaIX5/HJZs0syibNNZYPPNu0
vZ59hoLe6/1C9p5qMrItSMXkeJ2zcQ0/fnfR6dNhWfd0/Jw277QK/YT7j5ntNla9G2lqXKvS0jm0
couWO13T+UwtU5nvh0bUaoRs9YZKdN1pkq8Mgb+L20mLPX/bqrTbFhv+9pc0IP3nsGqNpnAIavWE
Ag+LT/PXOwgfo35IUBl5bEB/dRiFSIGoMJTPWklGP33D40Ci2zEwGJyAocoB1N5kWQTalscwF73S
65I1F9I1LuJdIp8EOMXK/6HsTrksXUegSQAx/+Z0TwrjM5lywyREzifOVLWGwazUeOUGXcewYzxw
yCptk1/US/60UM5tWPrD57/EJhA0lHR/YRY0QjCk9xd6Qy+as3+MimkoNbBo/MzDgtnZQAPcuEJj
Yy1tCOFf7hT+xpkWH+tFWqyfKYmbMBxBKQvds53XmQfcJc7W9gXIaFGcyU7ifhMmCMXklJuH4B6Q
etxefkT813o0RfBwaQ6FNuFtI/z1ajhZ8gm5KrmxZ4AGlU9f4kL9sFHf8boTpE2n74V5d+8v2MvP
6WkoWaxP3CGJ9XusxraRCJmA92JrbgUiGMQ7lh2MVtHZPWd/t09kfcsIg+I0NVjTAEGbxzYN2dum
SNjttwP7W5PbkKh4kZdQWxg+8/u/d+AQazAZZATipUSH1fx5/ec/oFvtB2FRHs876iz28widQ+T5
MRr+cRcSBrr7FqVY4t6+g9UWtIaLmwRwMpiHkHm3ViDHj4no5XTID7pUVRhVZGLgwlBApbfC1mN7
Gmw6GuemsKCvzKjTbd4euRmCXIOL78zFNDaMI4Vm5233lytfs7uDFLOEjrKkzhz5lnfy2CSkWRnL
DFmC7Yw1yrSch5Bgu6kC9ZcSA4t6wypGUVBIFU97wQRZH6fSKxm7z3U0L7coIa3ofXd5FdWq2OIv
YYsDtFJLgk0DDbC81M1sC14BbtVpTwv2g1m6Omyk+kLh5exnKpusI/FESKUn2RLtgAaW2f7oHOCQ
th2EPl7VZs7//5vvS3FDXpmyusogF3mE4r1EZR7qOfJyi2aDmPUQTxgs5DoWvsbIZ/zktbxMnFJ9
NbNb4kNd94guR/ovsaUovvRJQLuWZ4uNBYlzscnaG3BE/efIgjd8DYghd18mGTLhNSzJGa/Dl6qF
k72GtVq1Y3RzFKJNrdos7Ne/tJJohO+mz+wKmkPSDkTXkGhug7gUmGfp9PEmX5yMGGpXQct4JRVK
3SQ4r9zJIjmQrO5qIJ4xqITW6ktRJECjOdjkdn0d0avNaTS9SKHreCgts1iovQ7WZ5LeHzHeS/tc
xatpgGQntNNy+SlTx8sBVvKB8Djc6T9gMOvn9TZVwCaH03J8m8cujiIPyQhhccSLysKbgosy4cLr
vqJmeJZ5F07bgTVFFLqGmn3RCtge40RnFLEXcG8Za+pDVuMqNbGMFoTJtlkWQ6NNZBQ17oYorVk1
j7DKBMhxGfZWrAuAGfgXW5D+MZI6h1zqThG0Em3pX8uiZA57WKaIN9ynAYWWW6izwfglujVyMC4f
f1YDFMGdhnjpyAklFcTALXhOkx+Jgz+fOG0zzmcveAqZfE2s7UHnEpEnWIraqWoPdvktT8tmMehj
SqWNgVGJrfhqRvISGz/LRmI71/OLqVwxIqbUnbr8CErr5Ti4JufkxTil2OuxiRHu4LJl53qCgNM+
LZcuch6yzdAeoWwyPxMdKKzZE41Ddg15HOKS5/Z6BjpSeBiaGyVb1HPCi0N0oXfV9nL4ToevWLR1
B67jHil3Xj7qw7LH4kGG2ylw0cCkQ3T1zV6b79asQtQgsMxfw3ttBk418BPvMgoKeODagCHLP7rP
H2I8hoTR4VwIzW4v7Yn6yc7Wc9RWYbVqQ/+HgSvMNPWy5yzguDstb5Dy9WRXnx2vT3EFtPpESUFO
8idb5N3G3KTAUAVsO3FTMF6J9kcs7x2Obasx4ijbHlwBfznltBJE3scgTm8I1hFUVTcj0DyYe3aK
SfWTisZtekPm/jPuX/8qiAP/q/omyEO1jNtc0J90nCsGxibd2ePBh4KoWnfsJU5QQBRSJ8O0xmcN
qUOaYf3Z1YGJMKjB9sHhUZKAroNY/O69sBTZ/10ocWklXLqDU7v8a+d2HmuvIk2GC9Q1xJKTww7g
NgptFuOq6yj4ynr856KX0E/OWCHQt1CrUqC97CBkxBhQgsAfu/eoM2cQl4Y7JiWmE0fSV6p/yFoH
KbicL0knuHch4IX1Fx8yJjdqrg6BnAtMuVp4EKa73tvSuwUSdfAgaCPPkGYuIqrF1dEa0QGxlTnf
owmyt//rKOrXcixJkcTDMdrdxmL88qJvLw1R1vwpoKX5AiXrj6Pk7v+QobzY2wqezPqu8459Ocuv
31/ijt1iey4crwAayyeGPF3Eu/97ayzIIxCI68L21KxvNTS0IHj54KmXDx7cxNdZpY2Vx1tvSmVT
uQjcL4L9WXG4I312OUIjQmSEOPo3Y2hUS+A7UjmPkF6YJ09rZCgYo7l/W/lhLsqzJ+8gXwwOyRpb
op8DAZHgYYGFzYzh+HD9oV0zoeVU5QxQXKZfFQ9KARbJHXmAAY5a9Mul/cagDzk8kHjGhjSEgx5I
M6WChQgl2VILO/JtpWJheimuftFtdjZCp3aYGMks8pKIfUyBsS9HydLSxGL5Tp7g4OdfR4FcDD+X
RicY1CrEWq4eWznUS17CUXrvfm3HWSZdKuYOYgE7I96dIMtbo1j73qqCtBwVl7rU6CEMcFpv1N1G
vjEP5arPeSlF4kc76vkVnlXFRFlIns1CELsqxQjQPErhafzsl0M8YAsBtrQ2tJa63+dWS5wN/Bz4
i3vzu9Qr2yGklg/qwVd5bsuy07/M0JKB8ZnEOyK69ubaVHfjrZURY5Qe7ckxcKreuYSKs9B31sYa
xB4NM1LROFq+KJ0okNMEQ5zw6R4i8C+muXXSVEakzlUfniQdoJzXcsUX2EHSIUhlikd9PHYmLZqP
O16q2PfCUNJvP2xrEA0v0sy36ED1NQfyiMEUjf1/5rtDm1urDOQponbJ37h/1ulKQy8XYSGJfVjT
4YyBLiNIrc0R7YqetUeHxIgUnQ4+9mafG2AFtEwf+vdITZrqUbCzPmBzWKND8BETYhrY/5HJ3VEb
1MbD5TeaNBT+N9gUIgfh/YSOHAOd9+T0VPKFLA7r/mUg5kvocjBAlGTESkDlcG2Y1ZEvtIn00Rft
zfsxRCdcUwt1dBCL5pUZMGMei/YOGyn6WO5qt4SKbpI7/Q+F/MhDxFKll948FuE4Tn8EcSHyg2WJ
cZ97F8dHC3lVoQuQMELlZB/XKwlYhTHuBrUFYRV3dxIAeytqlXsauhoad89K2kzaCklze68Kc5T+
m46If/CtgRRTwt/QLTo+X9+KTaiAuDG3VPjLdlMZx8pl3P3h8wXcurJ0gsQmMg3gsWx8EAURFue7
A1G5pRiVENSa6SOz9lODwS0q7pttMoQLfc9ExEhqVvI+fufHoeRsS1fvF+w02Y/qdAWXNLq4z9y5
iQCMHg4qBIblv18ght0/mzLifhixpfni1F83FO88XmHRluyvt36XIpzeMGXXtADcRjbh59PHXvOQ
Zk8ztbStSQXxAIkKRfd2ktGlkjHY5tUg54zz7XRvMHzF5BYo+AtpLz9lwqDv8tt766jph0WOwkVt
sZq/eCwk5VX49rjBWo0iYJze23xheEqMxkBImVzZsIzBaClO9aUYY4/H2stmef7CPrTt1yejCfDF
ugBwZ92yRDL3VWSudHvDS01MxBqmhmfNz4pbllzIBDlLMkjncxlMYRSpW3GmXbroQfJdjTsNdwWK
TjyNpNlWUBV+FSgUpETBYgyDXwyGuHEQdHHgbdwyU467JWiwaJgY88oX+b/5KqdlZFjK0j9Rpi2m
lfRGnroyBT1n65n6/+n3yc/5jHDiQqiV6N5Exbt9UV04NfvSfU7yNOLXG/BqYKKNepjn++sK6u+O
StjiC4MTtE/eJe0DEPyMnsELthqQynCdZiEOv5tJLAC5eqhY0XWAlSe9u5G85TVrYZRpwTQcQ12G
YNqxUPioIIQJ9IUotce9eSFbfqT3pr8xORvYxluOCEE+UcYJhu4Wt6SHgfaHniT8Y2fvRMYevxGk
I5/Uf+nhlt2D7rUhPEf9KHnkduLODOYqgU9WqytfAN4MyB/4Lg3k+EtWxoTic6TUWGVQfw/hpqrj
SnqZvNNKLiIzdnqJIFtHDfF4nrbCsRHc1MQ9cIlZFIYKS/WCY/89uRNWC6Exqum0zWB2aAyT/aKM
gZX7auMqbBpz/EwaEGugsb9yWzlgNZZHo+Rh61NEXsxMYbhS5zVhKWmsQv0RU5Y2zILR0o5E6f1d
Dp1H2GYN+uhKZIUrI7B/bil2oBuL7HSofR4kf4oLazqPerOERh+aQpZ2FFVGBCeiCehCXIKem3qB
R1FYiW2c1tgqIoh+9Z3dpOVfYPMpmcCOIzYjImoA5GYU/mZGujT0IbbkNBU9/AyhFHS7OTmb/T69
Ee7lcOcy2lw+JFN6PDHZCW459VCplNmC7nZydrHxk//UgW0fEg2i5LhivjkqPN0NhogKTJ8FEfxM
Ekuo1Missr/wNp2i5jiXR8zPKgOsmTPut1QmdkVB552IhAF5pqSfF8QnALDuyQLQBy3YVlSsMQPh
qPc/22sMedk6Mlg0frs4MeGi094mmUiolCo0I2duxwe8T0FfsKaPAC/56NFiDMgxTOuwbH4NrruR
3GIE42BuhHQ28H/UaKqEV3JPMJJ6gnSZXbj9AY/pm6WbioRmHSKdYnks+0+09k9TdXaBCuD37YlF
olIGZPmlxuju1hg8hROgJCTIQ5mYAuYPexkZmbtLLBSbNVDtL9w+++ILICrzx9SGZ5PMWcJuDyzx
sz7Ab2f2/c3pNiG2oYKSUosypxnXgpzmjnNKdztv/I1cRmj0SEZpEUfXgpLXiys6V6YqxqozyUMH
+OctvxgbylkWog8dafn5f7H+5+XOorgNkt92+J1ivdfsNKUXygmvjXS+HWem5/RIj4gAv8NDzr79
unKrup5f+BevZ3nvTEGkS/dHUTpRXLWh8RadTuqYbn0dH0VE4v1Zbo2nbBZLNZxNgMgOJOJ+IGFd
mdAwirMtCbEl5ralQCMsO4GeQJOq2qnkVhiqzukKSk0RCkyvtqTu0Ris3OBnyH8dtuq7J135KpiY
6T7lBUCesy4JfAtufpys/jOxQzcXDc4eGlvwoyiBCYMH6Y15IJD0a1bW7f6UJFRCyQGbHZHypaCH
SE+4jROrs4cKLM5ECpzCgR9bxDydEgVh0YUeeWZQeI/xHPBt+Hf1zhbu1bfX2XMQj8UzzGp7YIeK
XXtrlIYaGCZOpc1fY2Vze6bhq1l+ODa4/GVfKzlxA7fCLzeh4nMl57M1VRZFTFY96PL2G/HF8VE2
HNhjFgDF26jZB4AtRnfNwhX95WNIS2wLtwiYqyCqKjLb06Cotp+JTsv/1Xakbcdd1pjCLuHEsZWC
jWA0laeQ3xBVoqI9DbMFTiYXlYHyWpZJY76zxIF8zURkyXPixIPIUEKqMtQaVy4pv+tXJmgpr3kK
mIp03PCyjtBu3c3LDW5JhjjnPbc+ZxIh+/LmRoqSgBMPoY/1pIRwly2BimF0AuaJBKOMrqMlhjJ6
A1c39+JlGu54q8/tJMPdl7lnOkfExTxb334YruBzKYpDoS++T5BU5jKHCTCtiXKvuA6wwHj4PKas
7JMi6CaaGdinBHqSqCOh7G0kH+8CXkU5dYxOXh/qKcUKONR6pZjnB/BvVLfGefy9Yd0Vl4ov2Bwm
bmZSx1I7aK3ym8g0xyIKjRtZ7OV5FJap+NOcJC3j3ciT6ETJ2aSdd8yLMi3SufaezrmHhjG8tPrt
Y/IfigOxqQ8dpPtvXuhf5pY1BZP0Gisk7VAeYqDhX4qiF6wQrM1EORd2JCdiJSy+1XHZz9vZNVT+
If8p4OFw+Db3O9Nb3h92ZudC6c/BfwjpVUhz/3lyCCKCceJ5auDqF6H9YNM6SUJL3S8r9ILiahRs
swfuSvmuBFpOI13ROE032BhDbScpTkyC4I0uetUT8kU1UV5u3E+no6f8cIGAqAw5qjYn4Kk4LJwg
IWFmeRlyg7gK4fNRLrKg1jWphs1pV5/cJRA8z5+cDRkqOp6eVbDoCTCG+CSL/VGSHrj0ZTErngZp
vw5/yglsnKvWvtJm6L9BofM0tOiTeCnfq7IKJ7AqDo9IT+ibvpn2ZRux2uJcpvc5/tSOZXYH17UA
WvjAyqpBOWbo6YuQx3Vjge0CewpclE2LIg5Nn7tNY3YJtqKsdNoEPmbqHo4bJv+ZpGVjf+kHSpoy
ls+gC9y9f238wQZzZ8y+/fGY74tmBHtL6GG5qQdYqrKPHuycUlSo2h5O9XzOIgV6DL9UF+qpkEIr
9YvFdydAKKKcg+I3Oltap2for2p+xVA4fRI6sQy7FakwWLMlQc9rzc4Qh6w5MOmu/V77SKLBFJoD
45P4/lRnKs34aw2d6LipAZY0w2aVUNKZKJ+tRr//B0da1ec8U3QjlxizZMQbV+s9CQ9XP561DLEp
2F881/DpIxnNm6x0SKH1gwmWKdjh3pWlAd4JD0VPK48WOAjzu0WyIvVoEY20UwhvNAByGoHhEgPU
ffhlGZG8+t1XHdTqNrrRXQJlxAAAOJRdi4Jkwjg2fcTReA9U4tZiGdNPUvCXfZh55Cm5+Nt32k3+
4rkByiyrIRTb1wKDM/fhIV1yb5lfKa1LBpIXlrAHqSEosN6zT1XNwhVuJeI+UJlPaw5OMkteEpRN
ghKmhyD4/57O4wvwdg==
`protect end_protected
