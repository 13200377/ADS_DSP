library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.filter_types.all;

package testBenchFilterIO is

constant numSamples : integer := 512;
constant test_input_I : int_arr(0 to numSamples-1)(sampleWidth-1 downto 0):= 
(		to_signed(116,sampleWidth),		to_signed(58,sampleWidth),		to_signed(0,sampleWidth),	to_signed(58,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(57,sampleWidth),		to_signed(0,sampleWidth),	to_signed(58,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(57,sampleWidth),		to_signed(0,sampleWidth),	to_signed(58,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(57,sampleWidth),		to_signed(0,sampleWidth),	to_signed(59,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(57,sampleWidth),		to_signed(0,sampleWidth),	to_signed(59,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(56,sampleWidth),		to_signed(0,sampleWidth),	to_signed(59,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(56,sampleWidth),		to_signed(0,sampleWidth),	to_signed(59,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(56,sampleWidth),		to_signed(0,sampleWidth),	to_signed(59,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(56,sampleWidth),		to_signed(0,sampleWidth),	to_signed(60,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(56,sampleWidth),		to_signed(0,sampleWidth),	to_signed(60,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(55,sampleWidth),		to_signed(0,sampleWidth),	to_signed(60,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(55,sampleWidth),		to_signed(0,sampleWidth),	to_signed(60,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(55,sampleWidth),		to_signed(0,sampleWidth),	to_signed(61,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(55,sampleWidth),		to_signed(0,sampleWidth),	to_signed(61,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(54,sampleWidth),		to_signed(0,sampleWidth),	to_signed(61,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(54,sampleWidth),		to_signed(0,sampleWidth),	to_signed(61,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(54,sampleWidth),		to_signed(0,sampleWidth),	to_signed(61,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(54,sampleWidth),		to_signed(0,sampleWidth),	to_signed(62,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(53,sampleWidth),		to_signed(0,sampleWidth),	to_signed(62,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(53,sampleWidth),		to_signed(0,sampleWidth),	to_signed(62,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(53,sampleWidth),		to_signed(0,sampleWidth),	to_signed(62,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(53,sampleWidth),		to_signed(0,sampleWidth),	to_signed(63,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(53,sampleWidth),		to_signed(0,sampleWidth),	to_signed(63,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(52,sampleWidth),		to_signed(0,sampleWidth),	to_signed(63,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(52,sampleWidth),		to_signed(0,sampleWidth),	to_signed(63,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(52,sampleWidth),		to_signed(0,sampleWidth),	to_signed(63,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(52,sampleWidth),		to_signed(0,sampleWidth),	to_signed(64,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(51,sampleWidth),		to_signed(0,sampleWidth),	to_signed(64,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(51,sampleWidth),		to_signed(0,sampleWidth),	to_signed(64,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(51,sampleWidth),		to_signed(0,sampleWidth),	to_signed(64,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(51,sampleWidth),		to_signed(0,sampleWidth),	to_signed(65,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(50,sampleWidth),		to_signed(0,sampleWidth),	to_signed(65,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(50,sampleWidth),		to_signed(0,sampleWidth),	to_signed(65,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(50,sampleWidth),		to_signed(0,sampleWidth),	to_signed(65,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(50,sampleWidth),		to_signed(0,sampleWidth),	to_signed(65,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(49,sampleWidth),		to_signed(0,sampleWidth),	to_signed(66,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(49,sampleWidth),		to_signed(0,sampleWidth),	to_signed(66,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(49,sampleWidth),		to_signed(0,sampleWidth),	to_signed(66,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(49,sampleWidth),		to_signed(0,sampleWidth),	to_signed(66,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(49,sampleWidth),		to_signed(0,sampleWidth),	to_signed(66,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(48,sampleWidth),		to_signed(0,sampleWidth),	to_signed(67,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(48,sampleWidth),		to_signed(0,sampleWidth),	to_signed(67,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(48,sampleWidth),		to_signed(0,sampleWidth),	to_signed(67,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(48,sampleWidth),		to_signed(0,sampleWidth),	to_signed(67,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(47,sampleWidth),		to_signed(0,sampleWidth),	to_signed(68,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(47,sampleWidth),		to_signed(0,sampleWidth),	to_signed(68,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(47,sampleWidth),		to_signed(0,sampleWidth),	to_signed(68,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(47,sampleWidth),		to_signed(0,sampleWidth),	to_signed(68,sampleWidth),
		to_signed(114,sampleWidth),		to_signed(46,sampleWidth),		to_signed(0,sampleWidth),	to_signed(68,sampleWidth),
		to_signed(114,sampleWidth),		to_signed(46,sampleWidth),		to_signed(0,sampleWidth),	to_signed(69,sampleWidth),
		to_signed(114,sampleWidth),		to_signed(46,sampleWidth),		to_signed(0,sampleWidth),	to_signed(69,sampleWidth),
		to_signed(114,sampleWidth),		to_signed(46,sampleWidth),		to_signed(0,sampleWidth),	to_signed(69,sampleWidth),
		to_signed(114,sampleWidth),		to_signed(45,sampleWidth),		to_signed(0,sampleWidth),	to_signed(69,sampleWidth),
		to_signed(114,sampleWidth),		to_signed(45,sampleWidth),		to_signed(0,sampleWidth),	to_signed(69,sampleWidth),
		to_signed(114,sampleWidth),		to_signed(45,sampleWidth),		to_signed(0,sampleWidth),	to_signed(70,sampleWidth),
		to_signed(114,sampleWidth),		to_signed(45,sampleWidth),		to_signed(0,sampleWidth),	to_signed(70,sampleWidth),
		to_signed(114,sampleWidth),		to_signed(44,sampleWidth),		to_signed(0,sampleWidth),	to_signed(70,sampleWidth),
		to_signed(114,sampleWidth),		to_signed(44,sampleWidth),		to_signed(0,sampleWidth),	to_signed(70,sampleWidth),
		to_signed(114,sampleWidth),		to_signed(44,sampleWidth),		to_signed(0,sampleWidth),	to_signed(70,sampleWidth),
		to_signed(114,sampleWidth),		to_signed(44,sampleWidth),		to_signed(1,sampleWidth),	to_signed(71,sampleWidth),
		to_signed(114,sampleWidth),		to_signed(43,sampleWidth),		to_signed(1,sampleWidth),	to_signed(71,sampleWidth),
		to_signed(114,sampleWidth),		to_signed(43,sampleWidth),		to_signed(1,sampleWidth),	to_signed(71,sampleWidth),
		to_signed(114,sampleWidth),		to_signed(43,sampleWidth),		to_signed(1,sampleWidth),	to_signed(71,sampleWidth),
		to_signed(113,sampleWidth),		to_signed(43,sampleWidth),		to_signed(1,sampleWidth),	to_signed(71,sampleWidth),
		to_signed(113,sampleWidth),		to_signed(42,sampleWidth),		to_signed(1,sampleWidth),	to_signed(72,sampleWidth),
		to_signed(113,sampleWidth),		to_signed(42,sampleWidth),		to_signed(1,sampleWidth),	to_signed(72,sampleWidth),
		to_signed(113,sampleWidth),		to_signed(42,sampleWidth),		to_signed(1,sampleWidth),	to_signed(72,sampleWidth),
		to_signed(113,sampleWidth),		to_signed(42,sampleWidth),		to_signed(1,sampleWidth),	to_signed(72,sampleWidth),
		to_signed(113,sampleWidth),		to_signed(42,sampleWidth),		to_signed(1,sampleWidth),	to_signed(72,sampleWidth),
		to_signed(113,sampleWidth),		to_signed(41,sampleWidth),		to_signed(1,sampleWidth),	to_signed(73,sampleWidth),
		to_signed(113,sampleWidth),		to_signed(41,sampleWidth),		to_signed(1,sampleWidth),	to_signed(73,sampleWidth),
		to_signed(113,sampleWidth),		to_signed(41,sampleWidth),		to_signed(1,sampleWidth),	to_signed(73,sampleWidth),
		to_signed(113,sampleWidth),		to_signed(41,sampleWidth),		to_signed(1,sampleWidth),	to_signed(73,sampleWidth),
		to_signed(113,sampleWidth),		to_signed(40,sampleWidth),		to_signed(1,sampleWidth),	to_signed(73,sampleWidth),
		to_signed(113,sampleWidth),		to_signed(40,sampleWidth),		to_signed(1,sampleWidth),	to_signed(74,sampleWidth),
		to_signed(112,sampleWidth),		to_signed(40,sampleWidth),		to_signed(1,sampleWidth),	to_signed(74,sampleWidth),
		to_signed(112,sampleWidth),		to_signed(40,sampleWidth),		to_signed(1,sampleWidth),	to_signed(74,sampleWidth),
		to_signed(112,sampleWidth),		to_signed(39,sampleWidth),		to_signed(1,sampleWidth),	to_signed(74,sampleWidth),
		to_signed(112,sampleWidth),		to_signed(39,sampleWidth),		to_signed(1,sampleWidth),	to_signed(74,sampleWidth),
		to_signed(112,sampleWidth),		to_signed(39,sampleWidth),		to_signed(1,sampleWidth),	to_signed(75,sampleWidth),
		to_signed(112,sampleWidth),		to_signed(39,sampleWidth),		to_signed(1,sampleWidth),	to_signed(75,sampleWidth),
		to_signed(112,sampleWidth),		to_signed(38,sampleWidth),		to_signed(1,sampleWidth),	to_signed(75,sampleWidth),
		to_signed(112,sampleWidth),		to_signed(38,sampleWidth),		to_signed(1,sampleWidth),	to_signed(75,sampleWidth),
		to_signed(112,sampleWidth),		to_signed(38,sampleWidth),		to_signed(1,sampleWidth),	to_signed(75,sampleWidth),
		to_signed(112,sampleWidth),		to_signed(38,sampleWidth),		to_signed(2,sampleWidth),	to_signed(76,sampleWidth),
		to_signed(111,sampleWidth),		to_signed(37,sampleWidth),		to_signed(2,sampleWidth),	to_signed(76,sampleWidth),
		to_signed(111,sampleWidth),		to_signed(37,sampleWidth),		to_signed(2,sampleWidth),	to_signed(76,sampleWidth),
		to_signed(111,sampleWidth),		to_signed(37,sampleWidth),		to_signed(2,sampleWidth),	to_signed(76,sampleWidth),
		to_signed(111,sampleWidth),		to_signed(37,sampleWidth),		to_signed(2,sampleWidth),	to_signed(76,sampleWidth),
		to_signed(111,sampleWidth),		to_signed(36,sampleWidth),		to_signed(2,sampleWidth),	to_signed(76,sampleWidth),
		to_signed(111,sampleWidth),		to_signed(36,sampleWidth),		to_signed(2,sampleWidth),	to_signed(77,sampleWidth),
		to_signed(111,sampleWidth),		to_signed(36,sampleWidth),		to_signed(2,sampleWidth),	to_signed(77,sampleWidth),
		to_signed(111,sampleWidth),		to_signed(36,sampleWidth),		to_signed(2,sampleWidth),	to_signed(77,sampleWidth),
		to_signed(111,sampleWidth),		to_signed(35,sampleWidth),		to_signed(2,sampleWidth),	to_signed(77,sampleWidth),
		to_signed(111,sampleWidth),		to_signed(35,sampleWidth),		to_signed(2,sampleWidth),	to_signed(77,sampleWidth),
		to_signed(110,sampleWidth),		to_signed(35,sampleWidth),		to_signed(2,sampleWidth),	to_signed(78,sampleWidth),
		to_signed(110,sampleWidth),		to_signed(35,sampleWidth),		to_signed(2,sampleWidth),	to_signed(78,sampleWidth),
		to_signed(110,sampleWidth),		to_signed(34,sampleWidth),		to_signed(2,sampleWidth),	to_signed(78,sampleWidth),
		to_signed(110,sampleWidth),		to_signed(34,sampleWidth),		to_signed(2,sampleWidth),	to_signed(78,sampleWidth),
		to_signed(110,sampleWidth),		to_signed(34,sampleWidth),		to_signed(2,sampleWidth),	to_signed(78,sampleWidth),
		to_signed(110,sampleWidth),		to_signed(34,sampleWidth),		to_signed(2,sampleWidth),	to_signed(78,sampleWidth),
		to_signed(110,sampleWidth),		to_signed(34,sampleWidth),		to_signed(2,sampleWidth),	to_signed(79,sampleWidth),
		to_signed(110,sampleWidth),		to_signed(33,sampleWidth),		to_signed(2,sampleWidth),	to_signed(79,sampleWidth),
		to_signed(109,sampleWidth),		to_signed(33,sampleWidth),		to_signed(3,sampleWidth),	to_signed(79,sampleWidth),
		to_signed(109,sampleWidth),		to_signed(33,sampleWidth),		to_signed(3,sampleWidth),	to_signed(79,sampleWidth),
		to_signed(109,sampleWidth),		to_signed(33,sampleWidth),		to_signed(3,sampleWidth),	to_signed(79,sampleWidth),
		to_signed(109,sampleWidth),		to_signed(32,sampleWidth),		to_signed(3,sampleWidth),	to_signed(80,sampleWidth),
		to_signed(109,sampleWidth),		to_signed(32,sampleWidth),		to_signed(3,sampleWidth),	to_signed(80,sampleWidth),
		to_signed(109,sampleWidth),		to_signed(32,sampleWidth),		to_signed(3,sampleWidth),	to_signed(80,sampleWidth),
		to_signed(109,sampleWidth),		to_signed(32,sampleWidth),		to_signed(3,sampleWidth),	to_signed(80,sampleWidth),
		to_signed(109,sampleWidth),		to_signed(31,sampleWidth),		to_signed(3,sampleWidth),	to_signed(80,sampleWidth),
		to_signed(108,sampleWidth),		to_signed(31,sampleWidth),		to_signed(3,sampleWidth),	to_signed(80,sampleWidth),
		to_signed(108,sampleWidth),		to_signed(31,sampleWidth),		to_signed(3,sampleWidth),	to_signed(81,sampleWidth),
		to_signed(108,sampleWidth),		to_signed(31,sampleWidth),		to_signed(3,sampleWidth),	to_signed(81,sampleWidth),
		to_signed(108,sampleWidth),		to_signed(30,sampleWidth),		to_signed(3,sampleWidth),	to_signed(81,sampleWidth),
		to_signed(108,sampleWidth),		to_signed(30,sampleWidth),		to_signed(3,sampleWidth),	to_signed(81,sampleWidth),
		to_signed(108,sampleWidth),		to_signed(30,sampleWidth),		to_signed(3,sampleWidth),	to_signed(81,sampleWidth),
		to_signed(108,sampleWidth),		to_signed(30,sampleWidth),		to_signed(3,sampleWidth),	to_signed(81,sampleWidth),
		to_signed(107,sampleWidth),		to_signed(29,sampleWidth),		to_signed(3,sampleWidth),	to_signed(82,sampleWidth),
		to_signed(107,sampleWidth),		to_signed(29,sampleWidth),		to_signed(3,sampleWidth),	to_signed(82,sampleWidth),
		to_signed(107,sampleWidth),		to_signed(29,sampleWidth),		to_signed(4,sampleWidth),	to_signed(82,sampleWidth),
		to_signed(107,sampleWidth),		to_signed(29,sampleWidth),		to_signed(4,sampleWidth),	to_signed(82,sampleWidth),
		to_signed(107,sampleWidth),		to_signed(28,sampleWidth),		to_signed(4,sampleWidth),	to_signed(82,sampleWidth),
		to_signed(107,sampleWidth),		to_signed(28,sampleWidth),		to_signed(4,sampleWidth),	to_signed(82,sampleWidth),
		to_signed(107,sampleWidth),		to_signed(28,sampleWidth),		to_signed(4,sampleWidth),	to_signed(83,sampleWidth),
		to_signed(106,sampleWidth),		to_signed(28,sampleWidth),		to_signed(4,sampleWidth),	to_signed(83,sampleWidth),
		to_signed(106,sampleWidth),		to_signed(27,sampleWidth),		to_signed(4,sampleWidth),	to_signed(83,sampleWidth),
		to_signed(106,sampleWidth),		to_signed(27,sampleWidth),		to_signed(4,sampleWidth),	to_signed(83,sampleWidth) );

constant test_input_Q : int_arr(0 to numSamples-1)(sampleWidth-1 downto 0):= 
(		to_signed(0,sampleWidth),		to_signed(58,sampleWidth),		to_signed(-1,sampleWidth),	to_signed(-59,sampleWidth),
		to_signed(0,sampleWidth),		to_signed(58,sampleWidth),		to_signed(-1,sampleWidth),	to_signed(-58,sampleWidth),
		to_signed(0,sampleWidth),		to_signed(58,sampleWidth),		to_signed(-1,sampleWidth),	to_signed(-58,sampleWidth),
		to_signed(1,sampleWidth),		to_signed(58,sampleWidth),		to_signed(-1,sampleWidth),	to_signed(-58,sampleWidth),
		to_signed(1,sampleWidth),		to_signed(58,sampleWidth),		to_signed(-1,sampleWidth),	to_signed(-58,sampleWidth),
		to_signed(1,sampleWidth),		to_signed(58,sampleWidth),		to_signed(-1,sampleWidth),	to_signed(-58,sampleWidth),
		to_signed(2,sampleWidth),		to_signed(59,sampleWidth),		to_signed(-1,sampleWidth),	to_signed(-58,sampleWidth),
		to_signed(2,sampleWidth),		to_signed(59,sampleWidth),		to_signed(-1,sampleWidth),	to_signed(-58,sampleWidth),
		to_signed(2,sampleWidth),		to_signed(59,sampleWidth),		to_signed(-1,sampleWidth),	to_signed(-57,sampleWidth),
		to_signed(3,sampleWidth),		to_signed(59,sampleWidth),		to_signed(-1,sampleWidth),	to_signed(-57,sampleWidth),
		to_signed(3,sampleWidth),		to_signed(59,sampleWidth),		to_signed(-1,sampleWidth),	to_signed(-57,sampleWidth),
		to_signed(4,sampleWidth),		to_signed(59,sampleWidth),		to_signed(-2,sampleWidth),	to_signed(-57,sampleWidth),
		to_signed(4,sampleWidth),		to_signed(59,sampleWidth),		to_signed(-2,sampleWidth),	to_signed(-57,sampleWidth),
		to_signed(4,sampleWidth),		to_signed(59,sampleWidth),		to_signed(-2,sampleWidth),	to_signed(-57,sampleWidth),
		to_signed(5,sampleWidth),		to_signed(60,sampleWidth),		to_signed(-2,sampleWidth),	to_signed(-57,sampleWidth),
		to_signed(5,sampleWidth),		to_signed(60,sampleWidth),		to_signed(-2,sampleWidth),	to_signed(-56,sampleWidth),
		to_signed(5,sampleWidth),		to_signed(60,sampleWidth),		to_signed(-2,sampleWidth),	to_signed(-56,sampleWidth),
		to_signed(6,sampleWidth),		to_signed(60,sampleWidth),		to_signed(-2,sampleWidth),	to_signed(-56,sampleWidth),
		to_signed(6,sampleWidth),		to_signed(60,sampleWidth),		to_signed(-2,sampleWidth),	to_signed(-56,sampleWidth),
		to_signed(6,sampleWidth),		to_signed(60,sampleWidth),		to_signed(-2,sampleWidth),	to_signed(-56,sampleWidth),
		to_signed(7,sampleWidth),		to_signed(60,sampleWidth),		to_signed(-2,sampleWidth),	to_signed(-56,sampleWidth),
		to_signed(7,sampleWidth),		to_signed(60,sampleWidth),		to_signed(-2,sampleWidth),	to_signed(-55,sampleWidth),
		to_signed(8,sampleWidth),		to_signed(61,sampleWidth),		to_signed(-3,sampleWidth),	to_signed(-55,sampleWidth),
		to_signed(8,sampleWidth),		to_signed(61,sampleWidth),		to_signed(-3,sampleWidth),	to_signed(-55,sampleWidth),
		to_signed(8,sampleWidth),		to_signed(61,sampleWidth),		to_signed(-3,sampleWidth),	to_signed(-55,sampleWidth),
		to_signed(9,sampleWidth),		to_signed(61,sampleWidth),		to_signed(-3,sampleWidth),	to_signed(-55,sampleWidth),
		to_signed(9,sampleWidth),		to_signed(61,sampleWidth),		to_signed(-3,sampleWidth),	to_signed(-55,sampleWidth),
		to_signed(9,sampleWidth),		to_signed(61,sampleWidth),		to_signed(-3,sampleWidth),	to_signed(-55,sampleWidth),
		to_signed(10,sampleWidth),		to_signed(61,sampleWidth),		to_signed(-3,sampleWidth),	to_signed(-54,sampleWidth),
		to_signed(10,sampleWidth),		to_signed(61,sampleWidth),		to_signed(-3,sampleWidth),	to_signed(-54,sampleWidth),
		to_signed(10,sampleWidth),		to_signed(61,sampleWidth),		to_signed(-3,sampleWidth),	to_signed(-54,sampleWidth),
		to_signed(11,sampleWidth),		to_signed(62,sampleWidth),		to_signed(-3,sampleWidth),	to_signed(-54,sampleWidth),
		to_signed(11,sampleWidth),		to_signed(62,sampleWidth),		to_signed(-3,sampleWidth),	to_signed(-54,sampleWidth),
		to_signed(12,sampleWidth),		to_signed(62,sampleWidth),		to_signed(-4,sampleWidth),	to_signed(-54,sampleWidth),
		to_signed(12,sampleWidth),		to_signed(62,sampleWidth),		to_signed(-4,sampleWidth),	to_signed(-53,sampleWidth),
		to_signed(12,sampleWidth),		to_signed(62,sampleWidth),		to_signed(-4,sampleWidth),	to_signed(-53,sampleWidth),
		to_signed(13,sampleWidth),		to_signed(62,sampleWidth),		to_signed(-4,sampleWidth),	to_signed(-53,sampleWidth),
		to_signed(13,sampleWidth),		to_signed(62,sampleWidth),		to_signed(-4,sampleWidth),	to_signed(-53,sampleWidth),
		to_signed(13,sampleWidth),		to_signed(62,sampleWidth),		to_signed(-4,sampleWidth),	to_signed(-53,sampleWidth),
		to_signed(14,sampleWidth),		to_signed(62,sampleWidth),		to_signed(-4,sampleWidth),	to_signed(-53,sampleWidth),
		to_signed(14,sampleWidth),		to_signed(62,sampleWidth),		to_signed(-4,sampleWidth),	to_signed(-52,sampleWidth),
		to_signed(14,sampleWidth),		to_signed(63,sampleWidth),		to_signed(-4,sampleWidth),	to_signed(-52,sampleWidth),
		to_signed(15,sampleWidth),		to_signed(63,sampleWidth),		to_signed(-4,sampleWidth),	to_signed(-52,sampleWidth),
		to_signed(15,sampleWidth),		to_signed(63,sampleWidth),		to_signed(-4,sampleWidth),	to_signed(-52,sampleWidth),
		to_signed(16,sampleWidth),		to_signed(63,sampleWidth),		to_signed(-5,sampleWidth),	to_signed(-52,sampleWidth),
		to_signed(16,sampleWidth),		to_signed(63,sampleWidth),		to_signed(-5,sampleWidth),	to_signed(-51,sampleWidth),
		to_signed(16,sampleWidth),		to_signed(63,sampleWidth),		to_signed(-5,sampleWidth),	to_signed(-51,sampleWidth),
		to_signed(17,sampleWidth),		to_signed(63,sampleWidth),		to_signed(-5,sampleWidth),	to_signed(-51,sampleWidth),
		to_signed(17,sampleWidth),		to_signed(63,sampleWidth),		to_signed(-5,sampleWidth),	to_signed(-51,sampleWidth),
		to_signed(17,sampleWidth),		to_signed(63,sampleWidth),		to_signed(-5,sampleWidth),	to_signed(-51,sampleWidth),
		to_signed(18,sampleWidth),		to_signed(63,sampleWidth),		to_signed(-5,sampleWidth),	to_signed(-51,sampleWidth),
		to_signed(18,sampleWidth),		to_signed(64,sampleWidth),		to_signed(-5,sampleWidth),	to_signed(-50,sampleWidth),
		to_signed(18,sampleWidth),		to_signed(64,sampleWidth),		to_signed(-5,sampleWidth),	to_signed(-50,sampleWidth),
		to_signed(19,sampleWidth),		to_signed(64,sampleWidth),		to_signed(-5,sampleWidth),	to_signed(-50,sampleWidth),
		to_signed(19,sampleWidth),		to_signed(64,sampleWidth),		to_signed(-5,sampleWidth),	to_signed(-50,sampleWidth),
		to_signed(19,sampleWidth),		to_signed(64,sampleWidth),		to_signed(-5,sampleWidth),	to_signed(-50,sampleWidth),
		to_signed(20,sampleWidth),		to_signed(64,sampleWidth),		to_signed(-6,sampleWidth),	to_signed(-49,sampleWidth),
		to_signed(20,sampleWidth),		to_signed(64,sampleWidth),		to_signed(-6,sampleWidth),	to_signed(-49,sampleWidth),
		to_signed(21,sampleWidth),		to_signed(64,sampleWidth),		to_signed(-6,sampleWidth),	to_signed(-49,sampleWidth),
		to_signed(21,sampleWidth),		to_signed(64,sampleWidth),		to_signed(-6,sampleWidth),	to_signed(-49,sampleWidth),
		to_signed(21,sampleWidth),		to_signed(64,sampleWidth),		to_signed(-6,sampleWidth),	to_signed(-49,sampleWidth),
		to_signed(22,sampleWidth),		to_signed(64,sampleWidth),		to_signed(-6,sampleWidth),	to_signed(-49,sampleWidth),
		to_signed(22,sampleWidth),		to_signed(64,sampleWidth),		to_signed(-6,sampleWidth),	to_signed(-48,sampleWidth),
		to_signed(22,sampleWidth),		to_signed(65,sampleWidth),		to_signed(-6,sampleWidth),	to_signed(-48,sampleWidth),
		to_signed(23,sampleWidth),		to_signed(65,sampleWidth),		to_signed(-6,sampleWidth),	to_signed(-48,sampleWidth),
		to_signed(23,sampleWidth),		to_signed(65,sampleWidth),		to_signed(-6,sampleWidth),	to_signed(-48,sampleWidth),
		to_signed(23,sampleWidth),		to_signed(65,sampleWidth),		to_signed(-6,sampleWidth),	to_signed(-48,sampleWidth),
		to_signed(24,sampleWidth),		to_signed(65,sampleWidth),		to_signed(-7,sampleWidth),	to_signed(-47,sampleWidth),
		to_signed(24,sampleWidth),		to_signed(65,sampleWidth),		to_signed(-7,sampleWidth),	to_signed(-47,sampleWidth),
		to_signed(24,sampleWidth),		to_signed(65,sampleWidth),		to_signed(-7,sampleWidth),	to_signed(-47,sampleWidth),
		to_signed(25,sampleWidth),		to_signed(65,sampleWidth),		to_signed(-7,sampleWidth),	to_signed(-47,sampleWidth),
		to_signed(25,sampleWidth),		to_signed(65,sampleWidth),		to_signed(-7,sampleWidth),	to_signed(-47,sampleWidth),
		to_signed(26,sampleWidth),		to_signed(65,sampleWidth),		to_signed(-7,sampleWidth),	to_signed(-46,sampleWidth),
		to_signed(26,sampleWidth),		to_signed(65,sampleWidth),		to_signed(-7,sampleWidth),	to_signed(-46,sampleWidth),
		to_signed(26,sampleWidth),		to_signed(65,sampleWidth),		to_signed(-7,sampleWidth),	to_signed(-46,sampleWidth),
		to_signed(27,sampleWidth),		to_signed(65,sampleWidth),		to_signed(-7,sampleWidth),	to_signed(-46,sampleWidth),
		to_signed(27,sampleWidth),		to_signed(65,sampleWidth),		to_signed(-7,sampleWidth),	to_signed(-46,sampleWidth),
		to_signed(27,sampleWidth),		to_signed(66,sampleWidth),		to_signed(-7,sampleWidth),	to_signed(-45,sampleWidth),
		to_signed(28,sampleWidth),		to_signed(66,sampleWidth),		to_signed(-7,sampleWidth),	to_signed(-45,sampleWidth),
		to_signed(28,sampleWidth),		to_signed(66,sampleWidth),		to_signed(-8,sampleWidth),	to_signed(-45,sampleWidth),
		to_signed(28,sampleWidth),		to_signed(66,sampleWidth),		to_signed(-8,sampleWidth),	to_signed(-45,sampleWidth),
		to_signed(29,sampleWidth),		to_signed(66,sampleWidth),		to_signed(-8,sampleWidth),	to_signed(-45,sampleWidth),
		to_signed(29,sampleWidth),		to_signed(66,sampleWidth),		to_signed(-8,sampleWidth),	to_signed(-44,sampleWidth),
		to_signed(29,sampleWidth),		to_signed(66,sampleWidth),		to_signed(-8,sampleWidth),	to_signed(-44,sampleWidth),
		to_signed(30,sampleWidth),		to_signed(66,sampleWidth),		to_signed(-8,sampleWidth),	to_signed(-44,sampleWidth),
		to_signed(30,sampleWidth),		to_signed(66,sampleWidth),		to_signed(-8,sampleWidth),	to_signed(-44,sampleWidth),
		to_signed(30,sampleWidth),		to_signed(66,sampleWidth),		to_signed(-8,sampleWidth),	to_signed(-44,sampleWidth),
		to_signed(31,sampleWidth),		to_signed(66,sampleWidth),		to_signed(-8,sampleWidth),	to_signed(-43,sampleWidth),
		to_signed(31,sampleWidth),		to_signed(66,sampleWidth),		to_signed(-8,sampleWidth),	to_signed(-43,sampleWidth),
		to_signed(32,sampleWidth),		to_signed(66,sampleWidth),		to_signed(-8,sampleWidth),	to_signed(-43,sampleWidth),
		to_signed(32,sampleWidth),		to_signed(66,sampleWidth),		to_signed(-8,sampleWidth),	to_signed(-43,sampleWidth),
		to_signed(32,sampleWidth),		to_signed(66,sampleWidth),		to_signed(-9,sampleWidth),	to_signed(-42,sampleWidth),
		to_signed(33,sampleWidth),		to_signed(66,sampleWidth),		to_signed(-9,sampleWidth),	to_signed(-42,sampleWidth),
		to_signed(33,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-9,sampleWidth),	to_signed(-42,sampleWidth),
		to_signed(33,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-9,sampleWidth),	to_signed(-42,sampleWidth),
		to_signed(34,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-9,sampleWidth),	to_signed(-42,sampleWidth),
		to_signed(34,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-9,sampleWidth),	to_signed(-41,sampleWidth),
		to_signed(34,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-9,sampleWidth),	to_signed(-41,sampleWidth),
		to_signed(35,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-9,sampleWidth),	to_signed(-41,sampleWidth),
		to_signed(35,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-9,sampleWidth),	to_signed(-41,sampleWidth),
		to_signed(35,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-9,sampleWidth),	to_signed(-41,sampleWidth),
		to_signed(36,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-9,sampleWidth),	to_signed(-40,sampleWidth),
		to_signed(36,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-9,sampleWidth),	to_signed(-40,sampleWidth),
		to_signed(36,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-9,sampleWidth),	to_signed(-40,sampleWidth),
		to_signed(37,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-10,sampleWidth),	to_signed(-40,sampleWidth),
		to_signed(37,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-10,sampleWidth),	to_signed(-39,sampleWidth),
		to_signed(37,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-10,sampleWidth),	to_signed(-39,sampleWidth),
		to_signed(38,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-10,sampleWidth),	to_signed(-39,sampleWidth),
		to_signed(38,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-10,sampleWidth),	to_signed(-39,sampleWidth),
		to_signed(38,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-10,sampleWidth),	to_signed(-38,sampleWidth),
		to_signed(39,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-10,sampleWidth),	to_signed(-38,sampleWidth),
		to_signed(39,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-10,sampleWidth),	to_signed(-38,sampleWidth),
		to_signed(39,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-10,sampleWidth),	to_signed(-38,sampleWidth),
		to_signed(40,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-10,sampleWidth),	to_signed(-38,sampleWidth),
		to_signed(40,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-10,sampleWidth),	to_signed(-37,sampleWidth),
		to_signed(40,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-10,sampleWidth),	to_signed(-37,sampleWidth),
		to_signed(41,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-10,sampleWidth),	to_signed(-37,sampleWidth),
		to_signed(41,sampleWidth),		to_signed(67,sampleWidth),		to_signed(-11,sampleWidth),	to_signed(-37,sampleWidth),
		to_signed(41,sampleWidth),		to_signed(68,sampleWidth),		to_signed(-11,sampleWidth),	to_signed(-36,sampleWidth),
		to_signed(42,sampleWidth),		to_signed(68,sampleWidth),		to_signed(-11,sampleWidth),	to_signed(-36,sampleWidth),
		to_signed(42,sampleWidth),		to_signed(68,sampleWidth),		to_signed(-11,sampleWidth),	to_signed(-36,sampleWidth),
		to_signed(42,sampleWidth),		to_signed(68,sampleWidth),		to_signed(-11,sampleWidth),	to_signed(-36,sampleWidth),
		to_signed(43,sampleWidth),		to_signed(68,sampleWidth),		to_signed(-11,sampleWidth),	to_signed(-35,sampleWidth),
		to_signed(43,sampleWidth),		to_signed(68,sampleWidth),		to_signed(-11,sampleWidth),	to_signed(-35,sampleWidth),
		to_signed(43,sampleWidth),		to_signed(68,sampleWidth),		to_signed(-11,sampleWidth),	to_signed(-35,sampleWidth),
		to_signed(44,sampleWidth),		to_signed(68,sampleWidth),		to_signed(-11,sampleWidth),	to_signed(-35,sampleWidth),
		to_signed(44,sampleWidth),		to_signed(68,sampleWidth),		to_signed(-11,sampleWidth),	to_signed(-35,sampleWidth),
		to_signed(44,sampleWidth),		to_signed(68,sampleWidth),		to_signed(-11,sampleWidth),	to_signed(-34,sampleWidth) );

constant I_filt : int_arr(0 to numSamples-1)(sampleWidth-1 downto 0):= 
(		to_signed(-14848,sampleWidth),		to_signed(0,sampleWidth),		to_signed(14592,sampleWidth),	to_signed(29696,sampleWidth),
		to_signed(14848,sampleWidth),		to_signed(0,sampleWidth),		to_signed(14848,sampleWidth),	to_signed(29696,sampleWidth),
		to_signed(-256,sampleWidth),		to_signed(0,sampleWidth),		to_signed(14592,sampleWidth),	to_signed(0,sampleWidth),
		to_signed(-14848,sampleWidth),		to_signed(0,sampleWidth),		to_signed(-29952,sampleWidth),	to_signed(-89088,sampleWidth),
		to_signed(-59392,sampleWidth),		to_signed(0,sampleWidth),		to_signed(-29440,sampleWidth),	to_signed(-59392,sampleWidth),
		to_signed(-29440,sampleWidth),		to_signed(0,sampleWidth),		to_signed(30208,sampleWidth),	to_signed(118784,sampleWidth),
		to_signed(88064,sampleWidth),		to_signed(0,sampleWidth),		to_signed(204032,sampleWidth),	to_signed(475136,sampleWidth),
		to_signed(281856,sampleWidth),		to_signed(0,sampleWidth),		to_signed(385280,sampleWidth),	to_signed(831488,sampleWidth),
		to_signed(446720,sampleWidth),		to_signed(0,sampleWidth),		to_signed(511232,sampleWidth),	to_signed(1009664,sampleWidth),
		to_signed(519424,sampleWidth),		to_signed(0,sampleWidth),		to_signed(528384,sampleWidth),	to_signed(1039360,sampleWidth),
		to_signed(512512,sampleWidth),		to_signed(0,sampleWidth),		to_signed(492288,sampleWidth),	to_signed(950272,sampleWidth),
		to_signed(479744,sampleWidth),		to_signed(0,sampleWidth),		to_signed(465152,sampleWidth),	to_signed(920576,sampleWidth),
		to_signed(467712,sampleWidth),		to_signed(0,sampleWidth),		to_signed(457728,sampleWidth),	to_signed(920576,sampleWidth),
		to_signed(483840,sampleWidth),		to_signed(0,sampleWidth),		to_signed(475648,sampleWidth),	to_signed(950272,sampleWidth),
		to_signed(484608,sampleWidth),		to_signed(0,sampleWidth),		to_signed(473088,sampleWidth),	to_signed(950272,sampleWidth),
		to_signed(502784,sampleWidth),		to_signed(0,sampleWidth),		to_signed(456704,sampleWidth),	to_signed(950272,sampleWidth),
		to_signed(489728,sampleWidth),		to_signed(0,sampleWidth),		to_signed(469504,sampleWidth),	to_signed(950272,sampleWidth),
		to_signed(506624,sampleWidth),		to_signed(0,sampleWidth),		to_signed(452608,sampleWidth),	to_signed(950272,sampleWidth),
		to_signed(493568,sampleWidth),		to_signed(0,sampleWidth),		to_signed(464384,sampleWidth),	to_signed(950272,sampleWidth),
		to_signed(511744,sampleWidth),		to_signed(0,sampleWidth),		to_signed(448512,sampleWidth),	to_signed(950272,sampleWidth),
		to_signed(497664,sampleWidth),		to_signed(0,sampleWidth),		to_signed(460544,sampleWidth),	to_signed(950272,sampleWidth),
		to_signed(515328,sampleWidth),		to_signed(0,sampleWidth),		to_signed(444416,sampleWidth),	to_signed(950272,sampleWidth),
		to_signed(501760,sampleWidth),		to_signed(0,sampleWidth),		to_signed(456192,sampleWidth),	to_signed(950272,sampleWidth),
		to_signed(514816,sampleWidth),		to_signed(0,sampleWidth),		to_signed(440576,sampleWidth),	to_signed(950272,sampleWidth),
		to_signed(506112,sampleWidth),		to_signed(0,sampleWidth),		to_signed(452096,sampleWidth),	to_signed(950016,sampleWidth),
		to_signed(519680,sampleWidth),		to_signed(0,sampleWidth),		to_signed(435456,sampleWidth),	to_signed(950272,sampleWidth),
		to_signed(509696,sampleWidth),		to_signed(0,sampleWidth),		to_signed(447744,sampleWidth),	to_signed(950272,sampleWidth),
		to_signed(524032,sampleWidth),		to_signed(0,sampleWidth),		to_signed(433408,sampleWidth),	to_signed(950016,sampleWidth),
		to_signed(515328,sampleWidth),		to_signed(0,sampleWidth),		to_signed(443648,sampleWidth),	to_signed(950784,sampleWidth),
		to_signed(528128,sampleWidth),		to_signed(0,sampleWidth),		to_signed(433408,sampleWidth),	to_signed(951040,sampleWidth),
		to_signed(515328,sampleWidth),		to_signed(0,sampleWidth),		to_signed(439296,sampleWidth),	to_signed(946176,sampleWidth),
		to_signed(532224,sampleWidth),		to_signed(0,sampleWidth),		to_signed(427776,sampleWidth),	to_signed(949248,sampleWidth),
		to_signed(517376,sampleWidth),		to_signed(0,sampleWidth),		to_signed(435200,sampleWidth),	to_signed(941568,sampleWidth),
		to_signed(536576,sampleWidth),		to_signed(0,sampleWidth),		to_signed(424192,sampleWidth),	to_signed(943104,sampleWidth),
		to_signed(522496,sampleWidth),		to_signed(0,sampleWidth),		to_signed(430848,sampleWidth),	to_signed(942080,sampleWidth),
		to_signed(540416,sampleWidth),		to_signed(0,sampleWidth),		to_signed(419840,sampleWidth),	to_signed(941312,sampleWidth),
		to_signed(526336,sampleWidth),		to_signed(0,sampleWidth),		to_signed(426752,sampleWidth),	to_signed(942336,sampleWidth),
		to_signed(545536,sampleWidth),		to_signed(0,sampleWidth),		to_signed(415744,sampleWidth),	to_signed(942336,sampleWidth),
		to_signed(530688,sampleWidth),		to_signed(0,sampleWidth),		to_signed(422656,sampleWidth),	to_signed(942080,sampleWidth),
		to_signed(549120,sampleWidth),		to_signed(0,sampleWidth),		to_signed(411648,sampleWidth),	to_signed(942080,sampleWidth),
		to_signed(534272,sampleWidth),		to_signed(0,sampleWidth),		to_signed(418304,sampleWidth),	to_signed(942080,sampleWidth),
		to_signed(548608,sampleWidth),		to_signed(0,sampleWidth),		to_signed(407552,sampleWidth),	to_signed(942080,sampleWidth),
		to_signed(539904,sampleWidth),		to_signed(0,sampleWidth),		to_signed(413440,sampleWidth),	to_signed(942080,sampleWidth),
		to_signed(553472,sampleWidth),		to_signed(0,sampleWidth),		to_signed(403456,sampleWidth),	to_signed(942080,sampleWidth),
		to_signed(539904,sampleWidth),		to_signed(0,sampleWidth),		to_signed(413952,sampleWidth),	to_signed(942080,sampleWidth),
		to_signed(557824,sampleWidth),		to_signed(0,sampleWidth),		to_signed(399360,sampleWidth),	to_signed(942080,sampleWidth),
		to_signed(541952,sampleWidth),		to_signed(0,sampleWidth),		to_signed(410368,sampleWidth),	to_signed(942080,sampleWidth),
		to_signed(561920,sampleWidth),		to_signed(0,sampleWidth),		to_signed(395264,sampleWidth),	to_signed(942080,sampleWidth),
		to_signed(547072,sampleWidth),		to_signed(0,sampleWidth),		to_signed(405248,sampleWidth),	to_signed(941824,sampleWidth),
		to_signed(565760,sampleWidth),		to_signed(0,sampleWidth),		to_signed(391168,sampleWidth),	to_signed(941824,sampleWidth),
		to_signed(550912,sampleWidth),		to_signed(0,sampleWidth),		to_signed(401408,sampleWidth),	to_signed(942080,sampleWidth),
		to_signed(570880,sampleWidth),		to_signed(0,sampleWidth),		to_signed(387072,sampleWidth),	to_signed(942848,sampleWidth),
		to_signed(555264,sampleWidth),		to_signed(0,sampleWidth),		to_signed(397056,sampleWidth),	to_signed(942592,sampleWidth),
		to_signed(574464,sampleWidth),		to_signed(0,sampleWidth),		to_signed(382976,sampleWidth),	to_signed(941056,sampleWidth),
		to_signed(558848,sampleWidth),		to_signed(0,sampleWidth),		to_signed(392960,sampleWidth),	to_signed(937984,sampleWidth),
		to_signed(573952,sampleWidth),		to_signed(0,sampleWidth),		to_signed(378880,sampleWidth),	to_signed(934912,sampleWidth),
		to_signed(564480,sampleWidth),		to_signed(0,sampleWidth),		to_signed(388608,sampleWidth),	to_signed(933376,sampleWidth),
		to_signed(578816,sampleWidth),		to_signed(0,sampleWidth),		to_signed(374784,sampleWidth),	to_signed(933120,sampleWidth),
		to_signed(564480,sampleWidth),		to_signed(256,sampleWidth),		to_signed(384512,sampleWidth),	to_signed(933888,sampleWidth),
		to_signed(582912,sampleWidth),		to_signed(0,sampleWidth),		to_signed(370688,sampleWidth),	to_signed(934144,sampleWidth),
		to_signed(566528,sampleWidth),		to_signed(256,sampleWidth),		to_signed(380160,sampleWidth),	to_signed(934144,sampleWidth),
		to_signed(587776,sampleWidth),		to_signed(256,sampleWidth),		to_signed(366592,sampleWidth),	to_signed(933888,sampleWidth),
		to_signed(571904,sampleWidth),		to_signed(-768,sampleWidth),		to_signed(376064,sampleWidth),	to_signed(933632,sampleWidth),
		to_signed(591360,sampleWidth),		to_signed(-512,sampleWidth),		to_signed(362496,sampleWidth),	to_signed(933888,sampleWidth),
		to_signed(575232,sampleWidth),		to_signed(2560,sampleWidth),		to_signed(371712,sampleWidth),	to_signed(933888,sampleWidth),
		to_signed(590848,sampleWidth),		to_signed(-256,sampleWidth),		to_signed(358400,sampleWidth),	to_signed(933632,sampleWidth),
		to_signed(580864,sampleWidth),		to_signed(8448,sampleWidth),		to_signed(367616,sampleWidth),	to_signed(934400,sampleWidth),
		to_signed(595712,sampleWidth),		to_signed(5632,sampleWidth),		to_signed(354304,sampleWidth),	to_signed(934656,sampleWidth),
		to_signed(580864,sampleWidth),		to_signed(8704,sampleWidth),		to_signed(363264,sampleWidth),	to_signed(929792,sampleWidth),
		to_signed(599808,sampleWidth),		to_signed(8960,sampleWidth),		to_signed(350464,sampleWidth),	to_signed(932864,sampleWidth),
		to_signed(582912,sampleWidth),		to_signed(7936,sampleWidth),		to_signed(359168,sampleWidth),	to_signed(925184,sampleWidth),
		to_signed(604672,sampleWidth),		to_signed(7936,sampleWidth),		to_signed(345344,sampleWidth),	to_signed(926720,sampleWidth),
		to_signed(588288,sampleWidth),		to_signed(8192,sampleWidth),		to_signed(354816,sampleWidth),	to_signed(925696,sampleWidth),
		to_signed(608256,sampleWidth),		to_signed(7936,sampleWidth),		to_signed(343296,sampleWidth),	to_signed(924928,sampleWidth),
		to_signed(591616,sampleWidth),		to_signed(8192,sampleWidth),		to_signed(350720,sampleWidth),	to_signed(925696,sampleWidth),
		to_signed(607744,sampleWidth),		to_signed(8192,sampleWidth),		to_signed(343296,sampleWidth),	to_signed(925952,sampleWidth),
		to_signed(597248,sampleWidth),		to_signed(8192,sampleWidth),		to_signed(346368,sampleWidth),	to_signed(925696,sampleWidth),
		to_signed(612608,sampleWidth),		to_signed(8192,sampleWidth),		to_signed(337664,sampleWidth),	to_signed(925440,sampleWidth),
		to_signed(597248,sampleWidth),		to_signed(8192,sampleWidth),		to_signed(342272,sampleWidth),	to_signed(926208,sampleWidth),
		to_signed(616704,sampleWidth),		to_signed(8192,sampleWidth),		to_signed(334080,sampleWidth),	to_signed(926464,sampleWidth),
		to_signed(599296,sampleWidth),		to_signed(8192,sampleWidth),		to_signed(337920,sampleWidth),	to_signed(921600,sampleWidth),
		to_signed(621568,sampleWidth),		to_signed(8192,sampleWidth),		to_signed(329728,sampleWidth),	to_signed(924672,sampleWidth),
		to_signed(604672,sampleWidth),		to_signed(8192,sampleWidth),		to_signed(333824,sampleWidth),	to_signed(916992,sampleWidth),
		to_signed(625152,sampleWidth),		to_signed(8192,sampleWidth),		to_signed(325632,sampleWidth),	to_signed(918528,sampleWidth),
		to_signed(608000,sampleWidth),		to_signed(8448,sampleWidth),		to_signed(329472,sampleWidth),	to_signed(917248,sampleWidth),
		to_signed(624640,sampleWidth),		to_signed(8448,sampleWidth),		to_signed(321536,sampleWidth),	to_signed(916736,sampleWidth),
		to_signed(613632,sampleWidth),		to_signed(8448,sampleWidth),		to_signed(325376,sampleWidth),	to_signed(917760,sampleWidth),
		to_signed(629504,sampleWidth),		to_signed(7680,sampleWidth),		to_signed(317440,sampleWidth),	to_signed(917504,sampleWidth),
		to_signed(613888,sampleWidth),		to_signed(7424,sampleWidth),		to_signed(321024,sampleWidth),	to_signed(918016,sampleWidth),
		to_signed(633600,sampleWidth),		to_signed(7936,sampleWidth),		to_signed(313344,sampleWidth),	to_signed(918272,sampleWidth),
		to_signed(615424,sampleWidth),		to_signed(10752,sampleWidth),		to_signed(316928,sampleWidth),	to_signed(913408,sampleWidth),
		to_signed(638464,sampleWidth),		to_signed(13824,sampleWidth),		to_signed(309248,sampleWidth),	to_signed(916480,sampleWidth),
		to_signed(622080,sampleWidth),		to_signed(16640,sampleWidth),		to_signed(312576,sampleWidth),	to_signed(908800,sampleWidth),
		to_signed(642048,sampleWidth),		to_signed(17152,sampleWidth),		to_signed(305152,sampleWidth),	to_signed(910336,sampleWidth),
		to_signed(621824,sampleWidth),		to_signed(16896,sampleWidth),		to_signed(308480,sampleWidth),	to_signed(909056,sampleWidth),
		to_signed(641280,sampleWidth),		to_signed(16128,sampleWidth),		to_signed(301056,sampleWidth),	to_signed(908544,sampleWidth),
		to_signed(623872,sampleWidth),		to_signed(16128,sampleWidth),		to_signed(304128,sampleWidth),	to_signed(909568,sampleWidth),
		to_signed(646912,sampleWidth),		to_signed(16128,sampleWidth),		to_signed(296960,sampleWidth),	to_signed(909312,sampleWidth),
		to_signed(629248,sampleWidth),		to_signed(16384,sampleWidth),		to_signed(300032,sampleWidth),	to_signed(909824,sampleWidth),
		to_signed(650752,sampleWidth),		to_signed(16384,sampleWidth),		to_signed(292864,sampleWidth),	to_signed(910080,sampleWidth),
		to_signed(632576,sampleWidth),		to_signed(16384,sampleWidth),		to_signed(295936,sampleWidth),	to_signed(905216,sampleWidth),
		to_signed(649728,sampleWidth),		to_signed(16384,sampleWidth),		to_signed(288768,sampleWidth),	to_signed(908288,sampleWidth),
		to_signed(638208,sampleWidth),		to_signed(16640,sampleWidth),		to_signed(291584,sampleWidth),	to_signed(900352,sampleWidth),
		to_signed(655360,sampleWidth),		to_signed(16384,sampleWidth),		to_signed(284672,sampleWidth),	to_signed(902144,sampleWidth),
		to_signed(638464,sampleWidth),		to_signed(16640,sampleWidth),		to_signed(286720,sampleWidth),	to_signed(901120,sampleWidth),
		to_signed(659200,sampleWidth),		to_signed(16640,sampleWidth),		to_signed(280576,sampleWidth),	to_signed(900096,sampleWidth),
		to_signed(640000,sampleWidth),		to_signed(15616,sampleWidth),		to_signed(287232,sampleWidth),	to_signed(901888,sampleWidth),
		to_signed(658432,sampleWidth),		to_signed(15872,sampleWidth),		to_signed(276480,sampleWidth),	to_signed(902144,sampleWidth),
		to_signed(646656,sampleWidth),		to_signed(18944,sampleWidth),		to_signed(283648,sampleWidth),	to_signed(897024,sampleWidth),
		to_signed(663296,sampleWidth),		to_signed(16128,sampleWidth),		to_signed(272384,sampleWidth),	to_signed(900096,sampleWidth),
		to_signed(646656,sampleWidth),		to_signed(24832,sampleWidth),		to_signed(278528,sampleWidth),	to_signed(892160,sampleWidth),
		to_signed(667392,sampleWidth),		to_signed(22016,sampleWidth),		to_signed(268288,sampleWidth),	to_signed(893952,sampleWidth),
		to_signed(648192,sampleWidth),		to_signed(25088,sampleWidth),		to_signed(274688,sampleWidth),	to_signed(892928,sampleWidth),
		to_signed(672256,sampleWidth),		to_signed(25344,sampleWidth),		to_signed(264192,sampleWidth),	to_signed(891904,sampleWidth),
		to_signed(654848,sampleWidth),		to_signed(24320,sampleWidth),		to_signed(270336,sampleWidth),	to_signed(893696,sampleWidth),
		to_signed(675840,sampleWidth),		to_signed(24320,sampleWidth),		to_signed(260096,sampleWidth),	to_signed(893952,sampleWidth),
		to_signed(654848,sampleWidth),		to_signed(24576,sampleWidth),		to_signed(266240,sampleWidth),	to_signed(888832,sampleWidth),
		to_signed(675072,sampleWidth),		to_signed(24320,sampleWidth),		to_signed(256000,sampleWidth),	to_signed(891904,sampleWidth),
		to_signed(656384,sampleWidth),		to_signed(24576,sampleWidth),		to_signed(261888,sampleWidth),	to_signed(883968,sampleWidth),
		to_signed(680704,sampleWidth),		to_signed(24576,sampleWidth),		to_signed(251904,sampleWidth),	to_signed(885504,sampleWidth),
		to_signed(663040,sampleWidth),		to_signed(24832,sampleWidth),		to_signed(257792,sampleWidth),	to_signed(884736,sampleWidth),
		to_signed(684544,sampleWidth),		to_signed(24832,sampleWidth),		to_signed(247808,sampleWidth),	to_signed(884736,sampleWidth),
		to_signed(663040,sampleWidth),		to_signed(24832,sampleWidth),		to_signed(253440,sampleWidth),	to_signed(885504,sampleWidth),
		to_signed(683520,sampleWidth),		to_signed(24064,sampleWidth),		to_signed(243712,sampleWidth),	to_signed(883968,sampleWidth),
		to_signed(664576,sampleWidth),		to_signed(23808,sampleWidth),		to_signed(249344,sampleWidth),	to_signed(880384,sampleWidth),
		to_signed(689152,sampleWidth),		to_signed(24320,sampleWidth),		to_signed(239616,sampleWidth),	to_signed(877568,sampleWidth),
		to_signed(671232,sampleWidth),		to_signed(27136,sampleWidth),		to_signed(244992,sampleWidth),	to_signed(876032,sampleWidth),
		to_signed(692992,sampleWidth),		to_signed(30208,sampleWidth),		to_signed(235520,sampleWidth),	to_signed(875520,sampleWidth) );

constant Q_filt : int_arr(0 to numSamples -1)(sampleWidth-1 downto 0):= 
(		to_signed(14848,sampleWidth),		to_signed(-256,sampleWidth),		to_signed(14848,sampleWidth),	to_signed(0,sampleWidth),
		to_signed(-15104,sampleWidth),		to_signed(-256,sampleWidth),		to_signed(14848,sampleWidth),	to_signed(0,sampleWidth),
		to_signed(0,sampleWidth),		to_signed(-256,sampleWidth),		to_signed(14848,sampleWidth),	to_signed(256,sampleWidth),
		to_signed(15360,sampleWidth),		to_signed(512,sampleWidth),		to_signed(-29696,sampleWidth),	to_signed(0,sampleWidth),
		to_signed(59392,sampleWidth),		to_signed(768,sampleWidth),		to_signed(-29696,sampleWidth),	to_signed(0,sampleWidth),
		to_signed(29952,sampleWidth),		to_signed(256,sampleWidth),		to_signed(29696,sampleWidth),	to_signed(256,sampleWidth),
		to_signed(-89088,sampleWidth),		to_signed(-2560,sampleWidth),		to_signed(208128,sampleWidth),	to_signed(-256,sampleWidth),
		to_signed(-287488,sampleWidth),		to_signed(-5632,sampleWidth),		to_signed(386304,sampleWidth),	to_signed(-512,sampleWidth),
		to_signed(-445696,sampleWidth),		to_signed(-8448,sampleWidth),		to_signed(519936,sampleWidth),	to_signed(4352,sampleWidth),
		to_signed(-523520,sampleWidth),		to_signed(-8960,sampleWidth),		to_signed(534016,sampleWidth),	to_signed(256,sampleWidth),
		to_signed(-504832,sampleWidth),		to_signed(-8960,sampleWidth),		to_signed(504320,sampleWidth),	to_signed(8448,sampleWidth),
		to_signed(-474624,sampleWidth),		to_signed(-7936,sampleWidth),		to_signed(475648,sampleWidth),	to_signed(8448,sampleWidth),
		to_signed(-461312,sampleWidth),		to_signed(-8192,sampleWidth),		to_signed(478720,sampleWidth),	to_signed(11776,sampleWidth),
		to_signed(-475648,sampleWidth),		to_signed(-8192,sampleWidth),		to_signed(496640,sampleWidth),	to_signed(15616,sampleWidth),
		to_signed(-473856,sampleWidth),		to_signed(-7424,sampleWidth),		to_signed(499200,sampleWidth),	to_signed(20480,sampleWidth),
		to_signed(-485376,sampleWidth),		to_signed(-7680,sampleWidth),		to_signed(484608,sampleWidth),	to_signed(17408,sampleWidth),
		to_signed(-467456,sampleWidth),		to_signed(-10752,sampleWidth),		to_signed(498944,sampleWidth),	to_signed(29440,sampleWidth),
		to_signed(-480768,sampleWidth),		to_signed(-7936,sampleWidth),		to_signed(482816,sampleWidth),	to_signed(23552,sampleWidth),
		to_signed(-467456,sampleWidth),		to_signed(-16640,sampleWidth),		to_signed(497664,sampleWidth),	to_signed(32512,sampleWidth),
		to_signed(-482048,sampleWidth),		to_signed(-13824,sampleWidth),		to_signed(484096,sampleWidth),	to_signed(33792,sampleWidth),
		to_signed(-465920,sampleWidth),		to_signed(-16896,sampleWidth),		to_signed(502016,sampleWidth),	to_signed(36352,sampleWidth),
		to_signed(-482304,sampleWidth),		to_signed(-17152,sampleWidth),		to_signed(489984,sampleWidth),	to_signed(39936,sampleWidth),
		to_signed(-459264,sampleWidth),		to_signed(-16384,sampleWidth),		to_signed(507648,sampleWidth),	to_signed(45568,sampleWidth),
		to_signed(-476416,sampleWidth),		to_signed(-16384,sampleWidth),		to_signed(492800,sampleWidth),	to_signed(41984,sampleWidth),
		to_signed(-459264,sampleWidth),		to_signed(-16640,sampleWidth),		to_signed(507392,sampleWidth),	to_signed(49408,sampleWidth),
		to_signed(-472832,sampleWidth),		to_signed(-15616,sampleWidth),		to_signed(491008,sampleWidth),	to_signed(48128,sampleWidth),
		to_signed(-457472,sampleWidth),		to_signed(-15616,sampleWidth),		to_signed(506112,sampleWidth),	to_signed(52480,sampleWidth),
		to_signed(-473856,sampleWidth),		to_signed(-16128,sampleWidth),		to_signed(492288,sampleWidth),	to_signed(58368,sampleWidth),
		to_signed(-451328,sampleWidth),		to_signed(-18944,sampleWidth),		to_signed(510464,sampleWidth),	to_signed(61440,sampleWidth),
		to_signed(-468224,sampleWidth),		to_signed(-22016,sampleWidth),		to_signed(498176,sampleWidth),	to_signed(64512,sampleWidth),
		to_signed(-450048,sampleWidth),		to_signed(-24832,sampleWidth),		to_signed(516096,sampleWidth),	to_signed(70400,sampleWidth),
		to_signed(-464384,sampleWidth),		to_signed(-25344,sampleWidth),		to_signed(500736,sampleWidth),	to_signed(66304,sampleWidth),
		to_signed(-451840,sampleWidth),		to_signed(-25344,sampleWidth),		to_signed(515840,sampleWidth),	to_signed(73728,sampleWidth),
		to_signed(-465408,sampleWidth),		to_signed(-24320,sampleWidth),		to_signed(499968,sampleWidth),	to_signed(73728,sampleWidth),
		to_signed(-449280,sampleWidth),		to_signed(-24576,sampleWidth),		to_signed(514560,sampleWidth),	to_signed(77056,sampleWidth),
		to_signed(-459776,sampleWidth),		to_signed(-24576,sampleWidth),		to_signed(499456,sampleWidth),	to_signed(81152,sampleWidth),
		to_signed(-442880,sampleWidth),		to_signed(-23808,sampleWidth),		to_signed(518912,sampleWidth),	to_signed(86016,sampleWidth),
		to_signed(-455936,sampleWidth),		to_signed(-24064,sampleWidth),		to_signed(500224,sampleWidth),	to_signed(82944,sampleWidth),
		to_signed(-442880,sampleWidth),		to_signed(-27136,sampleWidth),		to_signed(524288,sampleWidth),	to_signed(94976,sampleWidth),
		to_signed(-456960,sampleWidth),		to_signed(-24320,sampleWidth),		to_signed(506368,sampleWidth),	to_signed(89088,sampleWidth),
		to_signed(-441344,sampleWidth),		to_signed(-33024,sampleWidth),		to_signed(524288,sampleWidth),	to_signed(98048,sampleWidth),
		to_signed(-451328,sampleWidth),		to_signed(-30208,sampleWidth),		to_signed(508928,sampleWidth),	to_signed(99328,sampleWidth),
		to_signed(-434688,sampleWidth),		to_signed(-33280,sampleWidth),		to_signed(523776,sampleWidth),	to_signed(101888,sampleWidth),
		to_signed(-447488,sampleWidth),		to_signed(-33536,sampleWidth),		to_signed(508160,sampleWidth),	to_signed(105472,sampleWidth),
		to_signed(-434944,sampleWidth),		to_signed(-32768,sampleWidth),		to_signed(523264,sampleWidth),	to_signed(111104,sampleWidth),
		to_signed(-448512,sampleWidth),		to_signed(-32768,sampleWidth),		to_signed(507648,sampleWidth),	to_signed(107520,sampleWidth),
		to_signed(-432896,sampleWidth),		to_signed(-33024,sampleWidth),		to_signed(527360,sampleWidth),	to_signed(114944,sampleWidth),
		to_signed(-442880,sampleWidth),		to_signed(-32000,sampleWidth),		to_signed(508416,sampleWidth),	to_signed(113664,sampleWidth),
		to_signed(-427520,sampleWidth),		to_signed(-32000,sampleWidth),		to_signed(532736,sampleWidth),	to_signed(118016,sampleWidth),
		to_signed(-439040,sampleWidth),		to_signed(-32512,sampleWidth),		to_signed(514560,sampleWidth),	to_signed(123904,sampleWidth),
		to_signed(-424192,sampleWidth),		to_signed(-35328,sampleWidth),		to_signed(532736,sampleWidth),	to_signed(126976,sampleWidth),
		to_signed(-440064,sampleWidth),		to_signed(-38400,sampleWidth),		to_signed(517120,sampleWidth),	to_signed(130048,sampleWidth),
		to_signed(-418560,sampleWidth),		to_signed(-41216,sampleWidth),		to_signed(532224,sampleWidth),	to_signed(135936,sampleWidth),
		to_signed(-434432,sampleWidth),		to_signed(-41728,sampleWidth),		to_signed(516352,sampleWidth),	to_signed(131840,sampleWidth),
		to_signed(-418304,sampleWidth),		to_signed(-41472,sampleWidth),		to_signed(531712,sampleWidth),	to_signed(139008,sampleWidth),
		to_signed(-430592,sampleWidth),		to_signed(-40704,sampleWidth),		to_signed(515840,sampleWidth),	to_signed(139264,sampleWidth),
		to_signed(-416768,sampleWidth),		to_signed(-40960,sampleWidth),		to_signed(535808,sampleWidth),	to_signed(142848,sampleWidth),
		to_signed(-431360,sampleWidth),		to_signed(-40960,sampleWidth),		to_signed(516608,sampleWidth),	to_signed(146688,sampleWidth),
		to_signed(-410112,sampleWidth),		to_signed(-41216,sampleWidth),		to_signed(541184,sampleWidth),	to_signed(152064,sampleWidth),
		to_signed(-426496,sampleWidth),		to_signed(-40448,sampleWidth),		to_signed(522752,sampleWidth),	to_signed(148480,sampleWidth),
		to_signed(-410112,sampleWidth),		to_signed(-40192,sampleWidth),		to_signed(540928,sampleWidth),	to_signed(155904,sampleWidth),
		to_signed(-422400,sampleWidth),		to_signed(-40704,sampleWidth),		to_signed(525312,sampleWidth),	to_signed(154624,sampleWidth),
		to_signed(-408576,sampleWidth),		to_signed(-43520,sampleWidth),		to_signed(540672,sampleWidth),	to_signed(158976,sampleWidth),
		to_signed(-417536,sampleWidth),		to_signed(-46592,sampleWidth),		to_signed(524288,sampleWidth),	to_signed(164864,sampleWidth),
		to_signed(-401920,sampleWidth),		to_signed(-49408,sampleWidth),		to_signed(540928,sampleWidth),	to_signed(167936,sampleWidth),
		to_signed(-413952,sampleWidth),		to_signed(-49920,sampleWidth),		to_signed(524800,sampleWidth),	to_signed(171008,sampleWidth),
		to_signed(-402176,sampleWidth),		to_signed(-49920,sampleWidth),		to_signed(540160,sampleWidth),	to_signed(176896,sampleWidth),
		to_signed(-414720,sampleWidth),		to_signed(-48896,sampleWidth),		to_signed(523776,sampleWidth),	to_signed(172800,sampleWidth),
		to_signed(-400128,sampleWidth),		to_signed(-49152,sampleWidth),		to_signed(544256,sampleWidth),	to_signed(179968,sampleWidth),
		to_signed(-409088,sampleWidth),		to_signed(-49152,sampleWidth),		to_signed(524800,sampleWidth),	to_signed(180224,sampleWidth),
		to_signed(-394752,sampleWidth),		to_signed(-48384,sampleWidth),		to_signed(549632,sampleWidth),	to_signed(183808,sampleWidth),
		to_signed(-405248,sampleWidth),		to_signed(-48640,sampleWidth),		to_signed(530944,sampleWidth),	to_signed(187648,sampleWidth),
		to_signed(-391424,sampleWidth),		to_signed(-51712,sampleWidth),		to_signed(549376,sampleWidth),	to_signed(193024,sampleWidth),
		to_signed(-406016,sampleWidth),		to_signed(-48896,sampleWidth),		to_signed(533504,sampleWidth),	to_signed(189440,sampleWidth),
		to_signed(-385792,sampleWidth),		to_signed(-57600,sampleWidth),		to_signed(548864,sampleWidth),	to_signed(196864,sampleWidth),
		to_signed(-401152,sampleWidth),		to_signed(-54784,sampleWidth),		to_signed(532480,sampleWidth),	to_signed(195584,sampleWidth),
		to_signed(-385792,sampleWidth),		to_signed(-57856,sampleWidth),		to_signed(549376,sampleWidth),	to_signed(199936,sampleWidth),
		to_signed(-397056,sampleWidth),		to_signed(-58112,sampleWidth),		to_signed(532736,sampleWidth),	to_signed(205824,sampleWidth),
		to_signed(-383744,sampleWidth),		to_signed(-57344,sampleWidth),		to_signed(549376,sampleWidth),	to_signed(208896,sampleWidth),
		to_signed(-392192,sampleWidth),		to_signed(-57088,sampleWidth),		to_signed(532736,sampleWidth),	to_signed(211968,sampleWidth),
		to_signed(-378368,sampleWidth),		to_signed(-57600,sampleWidth),		to_signed(548608,sampleWidth),	to_signed(217856,sampleWidth),
		to_signed(-388608,sampleWidth),		to_signed(-57344,sampleWidth),		to_signed(531968,sampleWidth),	to_signed(213760,sampleWidth),
		to_signed(-375040,sampleWidth),		to_signed(-56576,sampleWidth),		to_signed(552704,sampleWidth),	to_signed(220928,sampleWidth),
		to_signed(-389120,sampleWidth),		to_signed(-56832,sampleWidth),		to_signed(532992,sampleWidth),	to_signed(221184,sampleWidth),
		to_signed(-369408,sampleWidth),		to_signed(-59904,sampleWidth),		to_signed(558080,sampleWidth),	to_signed(224768,sampleWidth),
		to_signed(-384256,sampleWidth),		to_signed(-57088,sampleWidth),		to_signed(539136,sampleWidth),	to_signed(228608,sampleWidth),
		to_signed(-369408,sampleWidth),		to_signed(-65792,sampleWidth),		to_signed(557824,sampleWidth),	to_signed(233984,sampleWidth),
		to_signed(-380160,sampleWidth),		to_signed(-62976,sampleWidth),		to_signed(541696,sampleWidth),	to_signed(230144,sampleWidth),
		to_signed(-367360,sampleWidth),		to_signed(-66048,sampleWidth),		to_signed(557312,sampleWidth),	to_signed(237824,sampleWidth),
		to_signed(-375296,sampleWidth),		to_signed(-66304,sampleWidth),		to_signed(540672,sampleWidth),	to_signed(237568,sampleWidth),
		to_signed(-362240,sampleWidth),		to_signed(-65536,sampleWidth),		to_signed(557568,sampleWidth),	to_signed(240896,sampleWidth),
		to_signed(-371712,sampleWidth),		to_signed(-65280,sampleWidth),		to_signed(540928,sampleWidth),	to_signed(244992,sampleWidth),
		to_signed(-358400,sampleWidth),		to_signed(-65792,sampleWidth),		to_signed(557824,sampleWidth),	to_signed(249856,sampleWidth),
		to_signed(-372224,sampleWidth),		to_signed(-65536,sampleWidth),		to_signed(540672,sampleWidth),	to_signed(246784,sampleWidth),
		to_signed(-354048,sampleWidth),		to_signed(-64768,sampleWidth),		to_signed(557824,sampleWidth),	to_signed(258816,sampleWidth),
		to_signed(-367360,sampleWidth),		to_signed(-65024,sampleWidth),		to_signed(540928,sampleWidth),	to_signed(252928,sampleWidth),
		to_signed(-350464,sampleWidth),		to_signed(-68096,sampleWidth),		to_signed(557056,sampleWidth),	to_signed(261888,sampleWidth),
		to_signed(-363008,sampleWidth),		to_signed(-65280,sampleWidth),		to_signed(540160,sampleWidth),	to_signed(263168,sampleWidth),
		to_signed(-344832,sampleWidth),		to_signed(-73984,sampleWidth),		to_signed(561152,sampleWidth),	to_signed(265728,sampleWidth),
		to_signed(-358912,sampleWidth),		to_signed(-71168,sampleWidth),		to_signed(541184,sampleWidth),	to_signed(269312,sampleWidth),
		to_signed(-344832,sampleWidth),		to_signed(-74240,sampleWidth),		to_signed(566528,sampleWidth),	to_signed(274944,sampleWidth),
		to_signed(-355072,sampleWidth),		to_signed(-74496,sampleWidth),		to_signed(547328,sampleWidth),	to_signed(271104,sampleWidth),
		to_signed(-342784,sampleWidth),		to_signed(-73472,sampleWidth),		to_signed(566272,sampleWidth),	to_signed(278528,sampleWidth),
		to_signed(-349952,sampleWidth),		to_signed(-73472,sampleWidth),		to_signed(549888,sampleWidth),	to_signed(278528,sampleWidth),
		to_signed(-337664,sampleWidth),		to_signed(-73984,sampleWidth),		to_signed(565760,sampleWidth),	to_signed(282112,sampleWidth),
		to_signed(-346368,sampleWidth),		to_signed(-73728,sampleWidth),		to_signed(548864,sampleWidth),	to_signed(285952,sampleWidth),
		to_signed(-333824,sampleWidth),		to_signed(-73984,sampleWidth),		to_signed(566016,sampleWidth),	to_signed(291328,sampleWidth),
		to_signed(-346880,sampleWidth),		to_signed(-73216,sampleWidth),		to_signed(549120,sampleWidth),	to_signed(287488,sampleWidth),
		to_signed(-329728,sampleWidth),		to_signed(-72960,sampleWidth),		to_signed(566016,sampleWidth),	to_signed(294912,sampleWidth),
		to_signed(-342016,sampleWidth),		to_signed(-73472,sampleWidth),		to_signed(548864,sampleWidth),	to_signed(294912,sampleWidth),
		to_signed(-325632,sampleWidth),		to_signed(-76288,sampleWidth),		to_signed(566016,sampleWidth),	to_signed(298496,sampleWidth),
		to_signed(-337664,sampleWidth),		to_signed(-79360,sampleWidth),		to_signed(548864,sampleWidth),	to_signed(302336,sampleWidth),
		to_signed(-321280,sampleWidth),		to_signed(-82176,sampleWidth),		to_signed(566016,sampleWidth),	to_signed(307712,sampleWidth),
		to_signed(-333568,sampleWidth),		to_signed(-82688,sampleWidth),		to_signed(548864,sampleWidth),	to_signed(303872,sampleWidth),
		to_signed(-317696,sampleWidth),		to_signed(-82432,sampleWidth),		to_signed(566016,sampleWidth),	to_signed(311296,sampleWidth),
		to_signed(-329472,sampleWidth),		to_signed(-81664,sampleWidth),		to_signed(548864,sampleWidth),	to_signed(311296,sampleWidth),
		to_signed(-312064,sampleWidth),		to_signed(-81920,sampleWidth),		to_signed(566016,sampleWidth),	to_signed(314880,sampleWidth),
		to_signed(-325120,sampleWidth),		to_signed(-81664,sampleWidth),		to_signed(548864,sampleWidth),	to_signed(318720,sampleWidth),
		to_signed(-312064,sampleWidth),		to_signed(-82176,sampleWidth),		to_signed(566272,sampleWidth),	to_signed(324096,sampleWidth),
		to_signed(-321024,sampleWidth),		to_signed(-82176,sampleWidth),		to_signed(549120,sampleWidth),	to_signed(320256,sampleWidth),
		to_signed(-310016,sampleWidth),		to_signed(-81152,sampleWidth),		to_signed(566272,sampleWidth),	to_signed(327680,sampleWidth),
		to_signed(-316672,sampleWidth),		to_signed(-81408,sampleWidth),		to_signed(548352,sampleWidth),	to_signed(327680,sampleWidth),
		to_signed(-304896,sampleWidth),		to_signed(-84480,sampleWidth),		to_signed(565504,sampleWidth),	to_signed(331264,sampleWidth),
		to_signed(-312576,sampleWidth),		to_signed(-81664,sampleWidth),		to_signed(549376,sampleWidth),	to_signed(335104,sampleWidth),
		to_signed(-301056,sampleWidth),		to_signed(-90368,sampleWidth),		to_signed(569600,sampleWidth),	to_signed(340480,sampleWidth),
		to_signed(-308224,sampleWidth),		to_signed(-87552,sampleWidth),		to_signed(555520,sampleWidth),	to_signed(336640,sampleWidth),
		to_signed(-296960,sampleWidth),		to_signed(-90624,sampleWidth),		to_signed(574976,sampleWidth),	to_signed(344064,sampleWidth),
		to_signed(-304384,sampleWidth),		to_signed(-90880,sampleWidth),		to_signed(558080,sampleWidth),	to_signed(344064,sampleWidth) );

end package;