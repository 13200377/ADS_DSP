-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
PzDCqhDY+pJY3Qc3heaUZ1enWMwcXcgstZG11BfYmFO/ZX56d5hHU1Sk/gcbo/kSZUyRB+pOU6+F
mqpXiBnwjL+PmZLMlrVn2poDIFiXfSdgKrIphATjRV07ZH4WYSh8HIb8rF7pI1ZXlo42YITg2I6B
2y6SLV8Z72PCougIu5RuYiwLP5dX3kVchgGoB71sDKB+9awxlg5r9RyMPoqlOd5WlsiUB6SDXvUJ
0FP0Zw9+A3VAr4hnsYzJoWp+TsMRrzoB37ct6rqDjnfk/8aY1ttQaHgJIAi8CfvWPVNpzBGYlx1W
is/YtdHxzgG2oq8FDuU1aLFRvOkdCYK6G1IzbA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23888)
`protect data_block
GenqP2MqA+LUxbwH2ue/IQMoDrAf+F62OwzOZxqtBCFNCdriZUjziM4eIZRfdg/XxOazadQAUhvk
DogfYBqnytazs2LoHaMoHutMEpWn6cIPOzwAGKJxntb1xQDC05DnVkRmj3t2t6DZgSUOa01puP7T
xmynzFdTW49yNLLgmKdCaJrSLAIbLsMSnKChThuRQ8MwlnUCyrxZFglx7tlDwRR0EZBw2pczRAKS
m02KgOyrVZuQSTb3ebwsyClvrcLDd1tbielBjNq1wjn5s3iBFqAarN8MfW+BWw76w6XeNV8K0g28
+9appPObM6i2G98cTBz1q6DDLmrrcyKRYiyK8OWxOchrhEfKLdgntKCOvPAZ5At4hSvAWpDf4kmt
qjMA67TfodSpo7nqiwmhtiUju3NRJM1LM+HdbYmRlLEkUy7fvRZJTQXbvoEfgp0+yYux8ZfHgD3A
4n+JkZdYyYnTyFiEWvQeE+DLp7RJTcJxL3JaKCOhxpK9shmvITr9FWn7gpj8zynSATt0XvtRNS/X
JF3RMex5ROb+tTIMpRXDeVf7EL6Tc2kftydqdiCIudog7fX0k1lFwa1NvwUxG3nq6RXGqRZwGIjA
B80GVKi9B4TlAlqezZRskSSp383d6ffG4ar947ZVfWG+2XOsAaWY7mWw1JYf+PD/int5fcNc2vPe
/Fc7V5LLVcEyicV2fC3YKBewjq74yfu+R2n8WbLrKAks8JfgCtL5bgk6rqXH//YuWNQZ+SO3Bc1i
7FfID4+ZTstRFS9F0i1fwyaqb2e2Ju6dHX/ZKiyrNZMHZPnKxbKIcvdC48oD5Xj0x1BrvUscOMW8
2DmJ98yEvjzEttCczbBYQx7FP79MUwOBNpNZQHFH5Zo95iBTFGHSjqZBQj7fmo+rVaD+hQd0zbYt
F8DxMQhST7vxh6j1MQE3bd+KeYhV2gE6myy8UKunTeYErM+D1BivG+Rt/QQmYvkwm5ruVOEh+Kr3
1whW/hp4r7EhR6GjxlIzsKCITqxqgvZnmMU/DkqSQg9TefxOuw0fq8OBJ5dmtsRdAeOFocnQJMdM
xRPLfRwZajCOVRU/TVjSwODuTVw3KnW3YmTDN5Gg4DCScsQ6xO/w58VoEdzMfm9zgKf70LyESBAe
EPl4moWGrayNVdNLoJxsRj6ndtws/6JKoilYXF5vian55U3EVpSlOT9+Z1HVGLvr1bwl6WlRIYKq
+tPvSlTSIABMyoVZtSqC4dbrqItEgVaTF3YhwU5VHXrFz+EgmwSltHs7EWu27atmQLXswTulXehJ
THh/7Lz9tqLEW4iv7TFUQzZNvmsw0kK82c3Gb8VmgxAPxdOgmTvBhgC7MVDzyewFx8IUsLAoQANO
BcIFutpOMr7W1bWAGGH+SYXuaNhz29VST7P1ZkIy0mpb8h3rWUKi9Wzsmp/UYaSENesprQ1cngbD
U5N033NWVEvE8WrW9LahVyfNyJXUtkkZjeZqJKKgk2Mid0T1eYO4YWzkFoCrX52tWg9fiUC0nloj
AKW7wuETYTfM0uN3Ldjv2XFgsH/ilLgR0Sp93JSVRs5inuq4o1Fxrfb9+vb6uu+mJehBnbO5nRR2
9E/ZYxN/UdryQMs0ne3jNGt0q7QuvjN5ySIdl2Fnki2R9r8RystXGHQ7dlErwrAUCq034TIiy1dA
CXzv/jdmTUBjxLmJJC0aDSzhfcLinJXNdcSoShCEfqjwcTHmzJKyQNKBKqCU5r3uWC2EnFfCrjGC
JkemHcxzJD419LXBGkNz91+iaahGWvZYO8/Ib0t3iu1pTiy//QxjNUR3BehcrZhRgBPJpW+0OLVu
7FrNKXRvTNzrZI/fP6BrW1Lcsrv0i5uzS9HcuyNqZZZSgY/ulY5g9YNZzqRjCnjV+KHsbvVjOnbz
Oa6XhQufvUtYIOfGzviwF2NyNCsajvXD6CbaIY+I46Y5nzNenfsbCqDGTM0l2T/QQACDGxUP8KBe
6j9lyFGza/IoPjmIopw6GarTBhi4w5E/ZGQyMj7N3s4wiSPjCV2IbNowv5jxIUXXbjHlfcNxHxzK
E8cE5oSs9wdSX/MDU1wW0nFBbsEXAkP9Dy+uTHC8L/qgr9RZ8hy/mmWVw348Ndr1s3gXWdI1I48c
ASbHhfvjxKZeH5i/s1zvYCOHWfr+A2mF3raLHhxbXB26PNXFRkkt6X4fGVIBKNCaa01MngaAk1IX
EgXpnyIoO6pysweFawlgXKZ1g9YvMdpszFR+B0QaXEboCBpsrAFQZGktPzqH5D19ZrBtZ9X/q3yl
W0GM/KvCunTP1uJ0fa7EX+WRDt7NAwttXMh/JM4P11qB47EeQTE9H75Wmq/s2rH5AwP1M7ljAF8q
yPVQrf7W6B4hgKxDWYaPBpN5WKdznurNxnUTIdyrhYx3tnmdXMpY2WKhd9ZXW8OOr0xGjiTU8Qdi
F4t+ftln2LS7MTW36FK5UXhgixBvl4HcPFD/kk3oZZHRuBdp6Wv49lOeOgwzC6u/Wmoca/tXpj4b
TJsYvw6ws10sTMwM+mpgl/BrWjNVn1WQWUdUcnEtlr5lmOE94MiMGsCiWzrV/WVV3wDaXuOY7/VM
5qw+yERnAvA5EuG0ecZHd/hOf5SwZHel1IReHXcnAckBxgs3egpidiR91dUv3q6s5cLXwnVuocKx
eyOtWWVOHkHka5sM64lQHjES09DRelssC8u512WyLgqJKzZGfDGIKUVImD9FiZB+RkWJI6ygfLOS
GFp8w1znlmWzhLlY2IDBWUSKYuqmKIkXnmrt0DHL7EIG3GG/Cwq/+DlBGTh0kN1vhESQa6kswFRv
23DkD0X0yLpRaVciTJg4u6P/vMRHWx35qNr8LRXDh2+XFT4erRdiDobV3zV9JJn4x28/nJUGUbSx
3qFN02V4k9TyN8ysvfP8MFADIlOo/zA/n6N3gPDnd3mB5LSCxam67+i8ykfz7yZjJ7LYt1z0VD5d
c0/8qYpDPgqc3sgFxCXLaTavZOgy6dpvVGMe4Kzpzfg95xFFo2/+v8zq5Tz6/linK/8ckofBvkHp
XYcxRWP+QrcXPr4yL7VzqQP8BEUU577Gd7/brv4jJ9R6NhXnCOkpGv2VKnQSfFrxLFpbF7s1Yhkr
mHrZox9hNJvGBzFFc9iopRkP5cXwqU38rokeJmhfBG6K2vIyo20Tgj901JgY65+7nM+b4FkpCfOw
vuSmFaEP43JeH0fnx0ZpQB2aV3VMd+HpepY5n6hN+CY6kJ47nYk4jhab6Zx97A123aFUC5rZiOMJ
YZG8bsFV0apB2xpvZG4CWtGSg9ueHg7H9g6tXFlmuoiJ2QcMINbimZyqQn4EBhGMVDDdmjAqvcy2
XZnfSk742N4/caqNKQeLJVj56biY2TRBrfKNp9yiq5yhVQRKDIgqin60greSK32zjuBvJidixkCg
yKGHF5owZZh4rlVjcOcd4hpNJZs8BWJH+jCM5H5bTaaC7B7Vk1BU3ZUrIpHu5OiW+OGpwjUtOMcF
IVjV92Tw0EpSY2wVCfBa/dHiCzx/Nu9aOWT8eEKLpopUl7UzvyioT+A7ET/UA8vVHs+JkgdkyEqw
HNF4BwNbNhUoOygWBsI26TW3qVmW3mNQFHsioVe8WKxewIzzjw2WzYfw67TunBemW+tV80IbfqxW
pPmtRrD1F9VT/jRTyKTUNOs+8CkkgMIL6mfcBpPnnTgDsYhRtSOobcgtw1gLI8dyGu67XxTuu5VC
9poTL3Od5fSOcXOle9oCjnJ0nPn3rENLooK1wcdznWEDGltcVXJN3XrBP7UU7id3jMl6QmUsvPVe
VOUqWQ172EeMJKNo6RXwYgVhPzTUOVncMY97AL9S6ZgJeGVjOj06Xi7yKPA4esoIdiVlies1lriW
6HUpoD5CFvcI0KGRQ1EMmMDj4MgMHXhVZanzdNffCNw/lCiUd6IfHcCaTvmX39qOF6SJkmWofWYD
gIcCuCt4u/9obGrfRDsMNQemhjif3IIWBBFophHw77VNvrXEtsQoloOeLcI2qRWD6JHKsb94VSay
AivXsSel7qE04N0XQrm6SE67myCQWOHhSGVR4KVw0vQwIBaftrxAz4dGfNS5F3WvHn73pie6JQHa
47QjPplxB4GqVDE0Ygcdwymq6jQbXNjO+b7Lrcy7tVYSvcVC9oRUQzECRKfHgVZ7fxDmSExTGT3S
vY2L4qO8Ig6ybsnMxH5oBoYY69O4Hpi1dbXZW3EaZKDEcSWwBeIAdGPGIHPIpR3q7BPujANprYtz
8OiEnvubSHMk0Rm6APt+kkXZONII+WZ9dkuLaYQHfrEdeGB3yPoUy+ijXrWyRgA71aczzskufvPy
ISXTZJpW57GhTU1jUuJZKobQ+ObUa4muvxLp9QoVASGEV0QJk9oytwSUsNBPzOVbZvBi4xBbEMMW
JQ22lFFU/lcLeu3/SqZiSvo/R09tLfrjZp7QBOFp+D6c/k5yUJF6opOnjxo5G8vKISgkAb2KN+pk
gWBUrAkA8tsxTqrA0LtkJiIk71mkOC6xWYGfx1Iko6kMJnsT8Yaze+HPyOWkBFk9LwCPpLsHRxYP
MCF/PbaHxwtToeu6InuoqeIdm/jPhx8emuKRQ78WbLgVlXQIbX6G2akRlWKRYcAXTxkG35rV7eom
wVPSvnR7kbenSP8IMgrS+pGByBfPN6sg64mXCBcTMe2pRyJUVqtcoJCReoaKbRGZkhZD/Fnl1iMr
BwvD7v3G1kn15Dn198Ii7ScidWYkCQOsFlMSBzCf9SonozpZ6eAJ9t3zWSxQ6qQiYIYj6sK537Y8
A/X/lz4JMHhfzF9168EqQOu9NOu3nDTyIHL0NqAqOpgI6x6OXSvOacI2ln5SN+muyOiVLt+UOJdZ
m/1G4/zep5L7lf/5DarDTrTyTU2XW5pkVHGrPx+jxdvwyoM2r8OBh5JWokNQCbAAD3o+1qE9wFfQ
ThDC37epNGfiOMwngis+NbkRXK3dAs0J3LQWC6YeaSbbYJpubvnN4ANw8Pb+Pqw/UoAMlw7EIstn
A4K/oD5TC+PwamvyTiKjv9vMHyRKceuKUdTV7sZNqNkof5FGmD9355lNxKE9oK0jJsV9214DfPod
qAT3bUaSAivGC+Mqrp1HDCIQPJAuyiHO6AYiqJqCXFdq0jpeJgMxqFGmqIXxqDuidGMSuzu5kaqe
n4JGtb4CsVc7/IZr1dsop++xhxT344XBq/l2CK1pLrilAU9t9LDITbDti6pb2YTbBvuf0cu3M19p
zKRFik/JgyzIKqaUStVFHGmBvx1QoIgMaXW9r11DKcHWV93Yt5hIxkHLNlgmxBo2VdJOIVCMVR/b
Of5+uHG4HVWJ0zfMrppWiXpiNVuTNF5ooWpKbB5uJWGc6QFxlLztkHrAbMKjxrtsS1H5uvvHYC5v
L0qy9JaDMjI8rMXcTX4e2MBXKmRiKw7GhwHbo+g95bs5cQ8gX7tNL68F5VxAWgQJNHe7GXlgyHTQ
siA322Y6VS/4UaEp3Y6k6cezSIw82n/abhFRcqmYxy51h6lt2/2Z3HnkPTgVHyDxfI7zlZCRFK7x
yEjtU40ciRjeptmZluajAghhhpgGRwjpH6KowKIeb//TUOcJ/AH3xgfyITh1mSDiET1sctw5256Q
MKQdNzdRe9WDXidV1wPzqXTR0SALlIDZTJmtb47GAXCbNbDpzfs7u7eLT0uikktuPGeu5OudelYY
ctTli/dVQh9bZiPclqi27Kwoq0nsnL3upBcgqhqXdhq82OaQEZDwKcBZ+40CSVBjdaOavI1TehMB
aRUQah4KM9jDfVa+2zRx/sIM0P8yjX5gGGHJPxUzJ1IuAmQFWu+7ddhAaORjRQ7qzQwlJwMtVWqz
xCIfP3K52SS6S9CRS8NEq8DApeagMr6Xc/q+Szj7XlR6cl9qTncPDE2O/PZ3kER3ZGjrS0OsWczg
axtGx5X1oHl3Gqd2J2rkfb/+FqaJ6VoLna+nBQSFbCVrXYl7SlxgzJy8JkWEXeShvArEZR08Vs02
2AC3Jf/TBAsCotUUJONok/goPZtNyWWzWUjfFxSKXcCD0keqJO6rqt1XeFpk4F0x53F/BzAVNuaN
pREQibnRuV7XMBiD/iOObqWmjEWHFAIhew/GutPjoPNjjH4dgZ3HluPKU1VaF1IQzKu0rrGaPAmj
2PVVj8zdtymlCqLtnNuaDGIaprbYmbB8WmiHuQ85w3JjypQz2Gdz1Cq2SWITvKed2GR+C4QPXAPs
BBfsP4WNji+e7BaqueACGb3xzw0WHKiGEvpbOPsgumUs32i+68+xf/AMRkRMK9DSFrCRYtqTxuX9
7bd30Ksd2xRODzNiT0Mee8+9qkLm1K7nxCgsue7uPHNqeNmkt1AZDPnAk0oCS1363W/GmUVlLhE/
7KtAeP2MLgK0VvebsnFGcJwBJmV7tkshKaUQ9Hi5uCrrjX0rcnAec3UyKDfa1w9RW3F7RE2kBgjk
71bsvyuEOzRik1EQEngee9XSIN7XujBFODq0kc65xTQzcC6/4FJHoqoXCljFZ/i+cUGwXnwCDlz4
kLaXWdfkmI19Y2JBZL0FO3UB690VQL29ftCA2vQHKPrP70lsTTXyG991rfU8QnObqtHbe/kSx6MS
2uKC+Oya9uwf5Ev2NT1omf1Et9K+QkaQz72r5mQdZ0hqbmV0Uu2EmN+lxRpH7/jJPPrKvS6xK0wc
WkYYSX1VHYjukdyl1Ku7AZmiCSZu48/6bQwrN9WdDDX0Agq/Ns0H7Ldcgr3bu8nCEXejMZzYMIMN
SblztC0deBQuC4hlUNwUnpl4khV3njH+ienEeKo+a/qg/XxN+WpNrz71IoKg9pL9nhPzwnT9fhYZ
IDuyP/09s2IUAwwCiVmpQGUAhHBA9n/oVV69vleS7I203y1DZnoTOMpHBq4Is+mJvYftK9ZPZbiL
BmcIMLZjj1iWgZUCPqNzVFxsjPTdlnNxABaght4fW0MzIFra6gvi/m/HoWCQcykxOWEj3fx5KPou
/RotxilrLBZZtHJju/5SNBFvC/+odoIzLYli5tevzBPtKygWLKz/wkvp0ZsGKUEuJUvepK0Njp1Y
ORrKfWvofza3gl+VfQwLCS7Oj8gdBvIHOrNEOLmNs67ELVgo25rdeXWy5eFjuMv8UfKea6LM5ZeW
zIZOkQ/YY/0NGzpCfcJZh6a4NBna5xkQLPdZXT9bTFtA1kblLRBHipTEXQ7o+6e7niqCIeypcbss
JzjhZpqaaWsUYJsUm8qYNgSOZWVuqrADRDK7LPpXQoaav7sidvz+QdesMWmb/clYg3gOSu8wp39D
3sIacKnDbnks6Ak73WH/IVwIZOTTaG7MTjDB/lZTZt4rXmXfPG4KbMDbfP3CgjEO3Jd926fYUbRO
xqgrsYm09oxOeqD3IQ9KE8dbhSU56Q6zNy09iacJw6CwVOZsX6ppahkR28iMwNgD44MXSq1vbFsB
x8A3J2s51vJET78uB1t05/SIB3q7IYbl8Y6W/Ta4mXWgac6RBfxUFCyp0BxjXKm7gGzr1A87W873
QKleVbI22wExSMaRKHjvx+LHqwspU9hFA6C8ZRbSzB+HuZ48OaOKsJ13Tme7KpfaxzfnX9IfmWFb
bgaqTv9mkxuHhncPEyMvMz/2za6W/1jptxjcRRcXqhnLYjyRWBVgl8fATacejq476ymmeJnL98+Z
xSKcu2AUDYITtrrdcx4PtSTLQLfOesjNbzCpP4E6HZPF8EF44BgaN03SZO1WJI3k/sk9DRyr0NVo
be8uvZiAB/HCoKNlgKC+c0kZSrgG/QhANWwqTGk4BplQn99MIazI6BIH73+Yxj+fPpsxYhgxeKOv
hpseG9mXcprQYheMTfEBbTxdAMPHHGb/K6ewyQsLnKcJpFCypyelXvsvce2Teakq2lvFcntohFSx
Y8kP/v8CZlXla8odxQZvxNbLXwn9UW/11i/YWdWtK/UNlnfr3bvfH83lC/nnOaHw6m8IZVi+H1Yb
p0oYrTYdC4ijOY+Xgc2Uta8U0b1fOxLE2vBP/jmKObKlX7IGeO6Zar/9xvqeqUE6Itawam6ByHpL
6RySoQ0KqJWGiToJlvdTnITjC+ihZl61blgoy+rnOBMcaxODbzbtG3CpN8Q0+3OReK4y1Bpj0DAk
KQPt6eXPn3dajiwcdE5qHOtC4eu2sp3uWJnaG2p4ivFdI7t6MKQ0aCieRN9ZKvbXAuf/Yct3u8Uy
4vieoXaJz/oQhgfXLHWcW+IkXfz+t7RH7j3wRh0Oti1uBpygCEEXPCQ7rs+qN6/y6XQtWA8TiDvp
kxVP6TPmiUop+CBahNVHZ2f1nGWBj/YU8GO1WfTrn8V8clUuIbUsQVtYdfJpRdDPQNqfrTFp2KTV
4vTOq/wJt5g8YpYD57jEQBGawA/r22C5G0Bp+No91d1Rcq3Pwf26SJ8zR+3VdeKeAOzqtUUFFA7O
gyrqTWBqhxpxuygLoNKu/93TbSL5HijWLHsTatQxQsz4A2PtgyBOOzsfq6MkBnVoVlvFuWfzn0gm
yMGTx39KfRbU+Ny41WItQlAOzTOwFgLObsPyip5iHQ1P5FvtXJzy9sBNfiMwOWSgZN2QDAU42xX9
n3Ug0jlXyWZ4SvY2U480KRrY19m5/kiqffCxO/XMw08yOJW4ECvQZnNAmHkfMEVLVImUVNbDcJOu
v7pS8trxtoe7rG0n4SIlwtGBGpAU7+Qa330M1imAQpdKPoSfbgAt09zcw1U2fDhqVPj4kHp6AtEE
+H3huQsZ7YGzfSoQsTaKPpodGLbWs21vPRmFpRtW97+J94YDC1ojbiFhBvK7m7HW0pK1sdqLw0d5
EIS6jxvq4DOoJQ1pvbGZUEp7GLPUubGhaRhXMVZ9t/X6hbx1jogXm9vukuVucIJAy5mUbdWO57CU
aNVxWSKzUC6sQ4u0diYSyKON949WdyaKdd5JifWjg8mSbiC7+5wi8VhOCNEumV8ffverJ0dpAjUb
eMWrjUUuteWf79nef0IrV0pjyi8NTleeALbbMROnpG+gPBZZJe7/smmyg927DoCftZt1nECNsUhY
ITZeJw6DU8GeaR8rd3ltmnRh14eyhxyi+TmUiGKvLhlip3TggT2eTGKTK+MM4/Jtm3PyBOiEjJKF
6Ltp86IYKJPC6mrGusF1eUg7+jo2nEZoQlLA2/LvYvmMhZZ+vmkE9BNUvuZxIHaeaBIKILDmpdvs
oDobcwUK/Qppz6pmvsTxNuYZ//4C7ofgn4JCVqXGcDXp5Di5CUb+VVfqAnrkDNWc1ChjyAtgj+no
XSUd1c3yxC+e4b9RRDC103HjssUTkjDswUlYhX6QrW3OorNZTcGdqNBD3nR1W8a7uVFO0r6+3zZi
N6g/euQ4RUZlVayI/iAb4E53FL55+GQ3FGzxFm7zraI07nbz+jOYo80QWOLZfOb7VenqgDDwdSqQ
qfF+Z5rQHfiiHYRWz51tpepvS9Yq3gql2TEqSh+8HjS/aqnFy4YevKK/3FwieRC4984hzkj/hDbh
x6Fhlgkr0q36abuL7wLtoIw/Zvq5VORxh7ukMPUn219y8075KrmK2dzA3tCtN15NAMd2+91mhy3e
NGglSP4yiLyXl3sc68KtC9hAEOeb94fuNYFQxNkLt/BvU6Qu8kfHBbeBVfc2VMEd8cxRU1qoqVSv
lDUTlU2z22bBnBDFz24MbCWOMdNKJ2AfIlyTpGyfzQEWVyKxUW2ZPOjq7u5n1kpdKftgxrC5xUIc
aXSbodyxRd0KN32kHFEWD6g3gsMxnh2rC0zL+0yB7ZITQZXQ7H1R10kOtRf1zACgY5gewfZZpyy1
piglyT0XOQStcRz2NBspSdmShpiSY1Souz1yZffMF7i2fb7hXj5pNkwBDmQUOwGGNYCHFEzTwYrr
hVonWd77LlNCC3kMstKbuWFw0mv6j11aGzSBHIxPbflvM1dg1VSLzBveqcr43O8rUv2ZAVQ6LK2m
jad02OXsbnYBsT6yz3DnyzMcAemqKPvjPuUvGfmEVhBRA8C9gaXHQQPITUvCYvrTn7HVLdDIOBpf
rsVYqsIfWNPlWOPBp6jmGvECU9ahSI2gzfhA0+7VMuriKpsM0D86nNiTlYXjYCMAXhxquh2ZCXBu
LCoKE/hqAq2dpfpLfBOPt9gO0N5c/I+JLNJ0lp7ApqDBiCarp/sUCWiHcs+W/OA4SrmzSKwvmUFE
Hdx3uJbgaiWy/mM3xs+cnUVOcbRnGbQ32hOUipB9OXJ148t5neURHRYHGbDoebhh3ZQpWgXAhmsS
XTELIELs26jPyCT2vHLBulg+dc2dGVJE3DXhmN99c+mQgCDnnlUnSFrlZ/lTdg3HeOB2LbgvVa8N
nPyNBrL3xmYVklj0ACRdVmbkROgBSnDZ2x5bzKZAtQo6OctB6PQgoRfnGB33G+r/zrRHUXrHo0uU
MDMjgz8qxNbR7ZCpcO3KDQujJdbeDn4DdQeEW2fKtBaZRijqr0WbG5vEeTWUeQWFewg74JH5N6fZ
6O1J6TTM15cdKe3VKZY6KX0GSpnMq0/CI1ZiXzvzDYqT2+BCDsOLb+Yhr2d9gofU4K5ZxTZqnMfd
OVmgwadS3FlTE3PtYkEZAINFNEONUEvUKYX1HNW8KezTVyHm3HajjYdwpTraDpTAHM5/QQGREWs+
V3mBd1aJIUxrcE+EzKkodW8hb5FLGPwAkULgfx1Ux6m+iYsjrpwjpAlSjp8+oL3KZZKtvo84AEmU
TttgLC/VE/iAJmx1etvLms0GrlVg7VaHcywlE1B1H9B+4Dax5n1tc3Rasf2ZP0rdiApL6DDOEUEJ
7/2E7cGyT0avIeBwiT9ZPHDJ7zCdLz0XtpeQzKdcgtOSiP6xuaGFNvuHRkMv1jtT2iemylZZS38Y
1TlGhN21u8NUV7FHQ9ew0SvJIkgbX5LKl2qby+BdUPPxVpJV014MWRsXhxfAKc4xdrklCy49bsqQ
WjR9fhsFXMyspOyTPUbr/R0OoA3ABMuMhXXqZesG4Cq0lk6kuEy4nQpl7x8c7M3mRzeOYeu3QWkL
ajAbvaNHxkIl8M6RQK84EpOsW/N0cvDSvbqihQss6z62+Zq6MBpDgQOl0eDvtziRwczHty+8Qljb
nImIjU70XUen7df3R+9Do6/4KlvnxvkhDl6lMAX/cDVMEDjxVVRVK6HIQqDoBLNT+TQ64nUgVEa1
2NRtexm+7jnr5WvwRk0/r/qbPY4VCfdA845zybkTNa9WCzyqUEvtr3CVd7NE6eCMMKBWLq5fCBH+
8r8Q+aeZpk5tF/X3j46r2ECkG8u5MYkbs11oeFvnruwk+yDBv1os231swF0+M2BL7sqki9/nxMx0
ArR91ULTqWwZvA2nJ3S6o+M9iAOVv3f6keTLqU41NNJgV2Iw9KThXYmymhq6XJztoEMxUt+Y5zYA
21zbTzkcTKG7ioY4xCbhnptkcnmfwh0O6cBIa3+NdbHqVOMj9RQepyR7CgD5DVhToNTRxTmcTFAC
oSBrfT6he11Z/PXznCMLsmTBV4Svyuto/uqTUjmLnytTSUKx4X2vQGSnyeusE6OUMj8dCGUGLDPj
ecFYqPO7fd3f7M1n/7GK8bCEUwrwgemrjDFuVzQIOAi9g3ecz7BCOOvvrhGWxLCalVk3wAGw/wMk
tfPhgz6hAwnDEM8nofkhAABtcgjL78Swm7D9o+/KlvlNEzrf8nePbQNWL+s1UzmX4b3bmCi3ML5M
dufCD+WZaiM0QcaoZkAqtgqw481/YGOtF4EbwJK1FG/RzKHphdDQ8b8TozVFCvsAb0UE07VP9jig
4xfauCxeefuGz/v3zrIAEGhJvCswjoAAj1Guy9LxIFBtZEoBpKam8Yl1DxDTY5a946/f4gUhNY1D
ztvzDF/k2OQIwDRkHXnFeHag5LOZYaLdUR6SR4NET4FHlmjs5NkBAYFVXVzrxq00YQohm4jB7Bqv
wXoO1/Kf198oN72h93EBcCq1Qb/o6tjfOk9q5k4aReNhUdhu76kpdetBQHF4LahGz/Owq4dASeEF
eiaLjHw2yF6eHSOkUhrV83AwcElOVvJHAcIOwgIltEnnIy6vvi8tRjAWLD1Xgl0oSyRre5UyESaF
ZH6hJj1eCr2j/XphPkE/x01nbe/nyC+euFDDW8FmJk7ALyj7ZWLNr6uylVgJBn6vGrUEYx+yokRt
/0+EdOaaHkk8KDi/DSJS3YpQJ00l9Erpm3mdR69N8qJGifUmFhAP4y16UOmgatik215qs3OXptpm
+pfzzA/FoocRcfMAl/NkP72HW5Q+RKbLZjl+CaAEELarBXqjXd577gUTtZwdrgqyiQbaNkH2rOyG
eSWr/Q7EBxX2ENZ8FMobc+4wCUgshfcSjEN6EU1lnUlJ4CbUfwwIaw0jH/TG+mpDZaWGeaH4Ipea
zrv7Hzknj66+wYnvrz+CocGY29G0sXkOT24fuu0MQo6QpOQIwTVpGK/xfxkuqXR5KkE869yQzh4l
4RcIfilViKlR6yEjpWrUnglJYb07hzFJrayUghpBSr7icA7QpG+FPaq+3znAzygbZcJJd0R2ol0x
iVV7bMQywYanpUxD718sb6hg5D0nKeiR5Df0gkgXrKuMzGIta0WPZAyR4hIwQG9AmcxbacdeoH6M
xh7BFu73yN3mDxsTzcfe1ATEoXXNR09fOPLiMoNZ6uDMyvrbbFArsVg5mli156Nkrr9hn19cSmPr
ZdE7E73nhHXeIEviAvljGlh/wCoBNrGb01WgnUGCX6F6WznxdiykzEJVGH3YP/KIXuuuufeOY0Qn
j5y+zH1DeRi0vruKhK7b6RjEuzZ+F+vLyJKvHbt8dENvy+P/doTL5AEMa6ZVUYTuEduDkOo6bGz0
r6Jf7+KcYty/9XiCGt8+KWy1t1CUBFZjNRX9skoeUKmJsx8KyFW6dchcdXA/Gxy8eimpQfqbRnRR
U5SIap+sCTX3L4l2RXBnST/dN0aFxDm9C6jt4cMWg9SlzYkw0v4Z3KysPvX1zn1ve6H3WkXomHPw
6coYG9g/1cB2Fh7ICY3M15UuhAufnSoQIqKSZ2KS2ZlisysDp8n1TvV1TbaexL8hHqk01z5JQrDw
ZZpivc4AlSpcXxQ+sxlrR6sHa3N9NVtIzH3b3GqHUwoyLjKg2yLYNJhpWXIiQoWKzNCEnhdG1OYU
OrwL4ids8o7U44ScXKXdBN+mxcPZhaQbOFdjVQq/lSIqn/FhUspAsGAy1ymGzRRxNSjrl4Stth6a
HUvhylF2HBVNdFU/8M02uViz27zZ3QEVa6fhqi/STbnDqTt4cUqzL44s8N31aXOppZQyO49Sfzw3
leYxUbPoeoaovuAadJlcdYak9yu6xPLMzABDgPH4cnx0AN6w40fE3Ei8AqqU7AQjyqT4SFTvfTD8
fKaBCp9NB0Pc2olXS2dNE0QKWkM4KiHkcFr2ubpvabx5/lH+9bmSYfDtOrOoGp2We3mTo44+bIKQ
8jMwMHI1W9zMJ0ba5jiWod9MVz+ZJJEz2sokEBDsYq0fObqZr+mRsKaRDwbuyLy0RO3wAE2g3oir
QYaQrgbICIw4gbkV2Gk+/FFPuYIpzc3ur3yvDao+minJWnjlhRTp/AxmEuwhnBRztNHnNYB43ZSD
CEIhgnpF9B4IRFKGppAOOa8otiZj0RmnHD7dQW/y+ZrPrvrauuFXe5w6g7152eLgAH5bUHWoQaVu
X5QSJ8deEGLN7ZV4VrTkJFKlL9VTJ8Og1lUjdm0O3xw81gCJz071DyNIm4rx+lVWz3Yk3KpP3nN5
NN1/UcEc80DiQY6N8QxOkAcH8ufNeNdbJIWzsXqze7A7xTfzgf961ACh/+FXzfAplus2jY1BUvI7
MWLTP53+j3DFDszXcooCbD2oQMJq28TREopu1+N4RtSFRSfBaXv4OYsumQdqmkYNKmFwwwWPMNy8
Dq4yuw1dK97l4d/GmW+fkLw8T2sFjekBXzhHEtaAyalq0YS1Y99w2eLR6lQiIo+BTH+vQgo55R+L
Y7950TV8Wm6h3jwsp/mr72eeY5tWE3FXPU6M4gUve1Vt4ePJfslavFU+onZx2x0D1vgF9ElKPaKI
8C4oCtZ49W8aCymB5eqYhDznLF3aL/Pgy29jAU1/J8faYJDCso5PduHFr+zrGYJrkY0hFbAAJytk
xZ0h2dcV9855NIU44HqczDlhgnqHsKNEHVejvh3ZlvxoMLnZaS8E9tSwHuyFpClgJowWRJgUW94E
bYNYhFLSRjGE917n3rs/WH6KHCS20udnfcL6N8Yj0nKwkC4oldss3qFpnQFAgh+37E0HFavS1oH/
YB8/dCm+OQh8BlzPTr0/xxicdAIQwMkCyzF+xL7al7eUnxFNpyZhh6kB1cgIza2Ms7GMwohYB86j
JdSKr8PJkP1s9o2s+DFD85GnbwE+D4L6zI8vHzmkJc+GlkP5RecxopWCFs/l/N5VykYsk2xtK4ee
mU7HhwPKfYEfsAYzN8OD+Kksb8T4+ZMcjPs2iqKUPqHPkNcvou/5QOkllYQg32f8r2KdJuCLDjN6
8C2lkxzTuj7Kp1EVAnnEyM9xGpSOdKgem+9ICwPWTRkvHj7XM0csUm7D5WtJ/0k+G4/8APfHxyX9
zXamstUtvGjCj8RFFl5RD8i9+HFlN6RfcSAxq5snDDEbe7Y6RVbcxqU6XKUmpvRaROZe8TEAwLhO
8qpi5gE9t9gDc/PO3gXukTA/p+jTp3ktK6dyIQcPynOBDCqPxcGfCdmrFYSBM5fPX5HMYiS6FocT
uCQy3+INr2IleO6wEdWwci7vixzAC+1IUubyhJDLdFWFO55DpFak2eSL6aroi3Hsy0WmxK+HbSgv
f0vW2URkX3cbcK6Y+4oqtlPgJZ4MdNmlidiR9WjV2U4B2J7Q1/7wFdb///4bXh8jn6T3/TSG89GB
+qO1NQ+NuSVXOTwoH9m7PWsJrxJReNbi/YtXxk9sKyauwAYvDcsvDKONJ4JQzcBnA9puqVQCVeC7
48o8FL39j97Shha1GnPDclEEUNfMumHuPK0X6yufoDYOcidxa/5EEauKZMKCxAHjY+cVdLU5WeT1
FQ6hFmBzT/FS46OTsR2YZNJUsqjiDRTnVqyERWnQv3GbiUWB3TN7BHc474UfU/loETBGl9ehd9pk
NyS+OmV7FQvH2LLVlgxyxR/3E8ClM2XL74uWRQQ8++RhUzLzTELsYckP8fbv1FR5ZG8GUtTJ3gde
u+LMs9kRm6qkSjG6SHTASYO5ZpLXCIvbZZD+PshCfy/F4xWH5Qfj9cJAtSdnbnLi7mayFSzAWBaw
1nzSc4PzmcEvpuxBOha8BuBCdETSE3qv0H80PkhCcOBaNHl8ApEeFLAT9r9FgrwSsyW7QYdgbelc
Lc/m4SEInOEciu4ZndX9O+zzAuUSBJEEWaS01SWj22XeIP4Sf/wR84TIAH/gXITNdTkMCkg0hxoi
tajYNglJXu0o6xc3yU7AOBW8awlNNQsnrxyzcUG35xw18uOiD04+vWkrV4wnmN01/F8UqTkbz7En
MUxIwwTspubrsGCQoxxTDut75/9dW1szN48GQp8rMDWv4mgyPBc1dIpRDQ1MXyop1WSArpn0CSkq
w95TrXPQv4ioAP0ONqAay0WXc3HCYstvsxFfGEIf45qEjIwlWrICXzlVMbdCcp+DUBBbxO/jWSdH
I3udEHiPS2UBClnIJNbHS8L9LvYThi8FrWSe3+nSvaNSkDUEgu83fMbCR4FVtX4GCrXpe82wqUFx
TE2uxGueuaQlM0KxRznggDm96FaElhWD1ajQT5Fuwkxzr1KkCK3/ERj76d1XEQjGrAfXD0lWrO9i
gOAfWWZUDGGzuIir0I6LRK1YiVP8T062MGW8QJ89YjxiIhN6sTzP+EvJAxJ2RU6qRT/roFtOfhdK
TFCPJRSBJvfayV7uUCDNiPOiStmE11UwIJ9DgMRYib03HmS5JS2nrnJtV2plc9AOlzue9ixaaX+q
P/5KLPJ6EDAWuRHszDZrHbeH1ZC2mD266TGnD333pHS8/3gvyRpTj44xKP6nMW7FfshkcJwe6tkC
EKvrPrIq4PKQhVw1m4RHHglkkR9Du+b6ogg5iGfU7x+VE+rkkkYXfZtv4PXt98dkpiI8asdP0aAf
ku/R5jhPle94pCRuw+4ZCQOZRJy0JBITj+7Ycn0d+Sumr+iJlBIjQ91m9W2jG9JTZc4sx3Ae5U2W
/1Toz73AQpKkMSuJFtpBdE7kmQ3jslisdVh8tOXCsJrg5vXKyjqT3KCEUbdqvxaZ2BbApmnROcFE
hhuRbKFJG+EXNydIuRzQmjUOMFQlZqmpcVjKiAHGJXsSCs7/N2ZNN13CCbgUYy5Y4LQetJvMcafZ
6lpykK5UC+yATV8cT8+Vbp2W8cyNhQ7P5sVpgU1/+sBCV59l6uNtAvXZdT1g1e2NurGV0VdYG0XW
f4LzhmTG8ovFc6lPtC5A07GISIRRPc1GNmMXFRe5Dhor7guVSMHqTGuNkVUyGTMSqPueno4vBLYF
YemuVCyU7Y2ar/SJH4YhjfkQD/2VlCowVd6WRVMGbs4agHXTYTI1jJMuu9LZiaB33C4WH9Shn/kI
wyX+Y4u1y5qwbbkfC7asEh8G6G9znreRNk5jUbnHtLbyzS1H0SB033Vibx2UndAnujdH6n5AvBIi
Wsjfj++rrVkK0L4nx5OHuu6rmvFnVr8Lge5dnTg0O17y4ttoPtFOAw+Aj6dMEYKLv15SZ0W7XdxH
egoKbxkjSEKHSTnfQwkdGJOb1A5GWtuhvjz42LHtea2tyywVIV75MCZI3XEyH/dHwnx6biLyFucB
s1Qvvj+YwFLHZSriuzT2dH/ABHmeWYMC5f9DDXwtFKQ9I1tvOkd2y/ZD4vWaSXCE7exeZzMRLTFi
l3AT/DTBSAliaOxJgV5C+RwiZwC0ZJcw0gQIgDdrHaltXIYFqd5P4dsarBJMmhCgs139Z2eNu2Un
k8AdHPN/ZeGTh2vl5uOlVUG9tuMQHBjQEklgohih9MO3D8+LZ0ggyH4/KVnWgLaFO0b35mN6qR7W
vCd9mRBjud4aFVlb8h6AII1RB5lYwW5Fu4KuTE3j/6rs40zImubaXb7iEqpm6jGzlLv3Ds03vag9
/B93fcTrujzpZfqn+mlJaEL7KIIE13iJhdaEJUtnKQuGvjTWKhi54LpSEWoe00Jag1HTep3S4osU
C7OyibVDSW/7cJi5t8DVnCx6dyurDqZ5jZKwnZxSc5GSZTLRTSozzHj1ZvOcPPihf8Y3HTZ4MPna
rbhAvqNP3B20LVi7QN+5zhyAGyBk/nilNKzhHs0Uo1UPtR4yW+gNLYkHkFOE2uBHxoGT6LSkyc+3
Qwr4PRv3FrTUtG6caSA4wG0pvVh/mTX3w2qbdaiH82tfFFg/GGhcTVTrzkJq5CALMyIclPSC5tzK
J7JHErlynmQWVIJeSB4XTRgCmBrXZMdVmlFq8Y9c42P6FFuCxjljCY10CE4Dda2FEjrM36ZEqU3N
HaMICnVWHh5eRqI3B0NZsJtj6fDRmbaHDaBA1LYFIRlfPqc5B5uGunQjZwitGwZgPZtYuxL6Sp1G
sf7sBprydxUpTAAFZVHGYxk9Xt4ls0CIbwq4HTzQoy8HS959ogCO0XEZpYfTW46IA+Nj1XblH7yE
jbceqVUf4JkbCcUgzR117YWBH9LknLUFE49AlbR2f1ScoH6YER9mCfpXZ4kVZVmcQAW2rE4e5SGG
aBEeMD3oYqG/GlFmSVOM1DTBb7hmGZsSPCs12rgdi+Es9/xdS7wwhnSHxDMKqdg4Ir5wHGGoeZke
kr8ZU+VqDXqD3oXqlIsb1xFdcHDrdMvFCsoOJyomP3rvNCIRqa3LJ1xWGQcIhCM9u/OjjDmBXVs9
IZ0Oro9QFnEbEiHRD0J1Awp7Kv/aZx5mbipLv+bqezMDdcRuZJoTxwVlTRre6/HTcaUuMwwhG9HW
0/rgQdXyeJdeTvsny4A+SDactZlcryJekfhNV13Ri87fsQ45B7C8jC1WBwwzxm0y4h3g8APV581K
pmySHe/BWaC0uqCdMT9e3PBRNN+jNpZ4CAJoVzytVTPLWGm3/y9Y1QRSMSCpsdzTIY1WZsxlszxn
LNg72oFM+/mkCIT75azYJ3fsKeZtJe6Vn1HVDpXR6OkmcNZCcuOoeJt4+GhdLoYNkIMS9jg0Q91e
/EOLKoS5N/2j7Dnf1IN4SoUKvKeJ1IeZdeuuI1ypvGyVkOqQsFumKSqQEK/s87HXAe7er1QyTqXk
yUfGcjhiZsoH4MGoKcz1lSbZPSt892yVH9DSCeDJSMlgStUq8wv0Y1fpRvYb8GDcHFKdyh+axLXy
U8OXadJjSlZTgMhKyaGGnZ7q0pyH6aiZ50CerlOncjoRdlgVDsiAmNrp5UP9UM1RMjm+nLCJBTN5
S8fXoziNRe/E1Dm+mzcRzb79gvVtG8QPNc8G7rBAvZ5fXDW+culcMoarwWlCoNHLIdopApZzqj5k
CYYYVeqHP7WTMOqLZd4PH1S9JFYV1ZTX8GecVBADiKcVNeNuCPAhHQU5wkK5KiEaFunxaMCUBwTG
PbBRPeaVLVD4DpH06Bw4HC0o7vkfA7nIAFTwKO0khcHxS/+WnKgPv4vSRsZjNWSH2EBzJf1ccJ2G
0RGgbk3xhRS3Rx70kPAVEP8tCLdIgXXypejwdUTPZsTBP1wn1R9VWH9YGXMV72oHTjLcQojC4Vkr
kV2W3kffLsWyxzweLdGyPopH/mHjUCRpN39aOhxYGa96vgpitAy/v/b1KyVASReHr2g0t66NfwYr
DkNNeVfHM4ls+JlAMmHa+Syo9w8tIxsDnX6SA/sy+IeSTJd4LMvgiS9hlHY/TeBlJOF03+2UOa9n
gtAedJ1wPiy71FRpIOQlnZStpSEkGQ+lxZJU187F0PjCdxKVGuxWxLSqWqxX1cG3kodXaOAnmkz7
24/WYlNLwBiksvuSlE2DpLgftTYje42YEc9Mm1LgPMJekKwXbevozccRaf3aOtqaTsOAX5EJrjvC
+YPxJGq2F0HYByc2NLdiPB72bogei4AXWpSwy4i1j/6dOi+Nd0vwLSJhf6O9EVYcDU7W4RYEK62L
8FobDf6siXW12fxp8ZqjMa2uRzeDzLviPD/1fbNKArvaJB5c859ATedravzj0EWSGL78heuXhUki
1DAMbBOv5za1wyZt0DIKjKD0f29sCQRqhOw4FWhAuljuOXdE6gk+hCAOUza/OVMg6mdbQShdsbZB
hcI76Ur1wU9+kNQqy4Ut4xM1stp24qIZvqRbPUbhLp+nH8TgXHG7u3cN6tqOCqmLtixQbVd/JgYW
KAcdR6ld+Rl820KdaRfXz9C5OLLT4Gk7ZVoCuss87bTRAlO4OtI3cvNtDUj/Fc/Vg3jd4AMc82dD
ZrwEPjqxxl6EneKb53mo2iwhij3mFcKv1mPCVuX/4Umb3cSghzH5FXUf0wA0BueawRWtZEyfpyCM
tfFgZ+zp9Cq71nH3ywo9ecAAzEE7Qkp/o4elpYszaRMeDGKThSlD04Ed7WbXs1CN9uU4dx+MOZju
iyVm5tcSRIXID2YCglTf9VBIv0YO71N8pYDuWSUZx1TtQLuojEvJG1Gvsl6vCA43RsJAE0m7KEt5
d6DaqFtgdUFnv/oCK5kC7CQD3MRpvovIenEXuKo+KQPqHEKsf5WMUa3MMRvVf4TdbnuabKN0yDKB
37FkcufooAbraNdai65XG86IFW5QifVKI8ek5jNHMG1YFYp8spnmisc7Hgd2wU3mKH8VTsdg44hd
LDRa/jwudYIPscM5c6Gc7YdiV5U//4Fas+Ej1tBQjtJg1i0+/Vinbyw3MMPKYjyHLLeXkco0a2Kh
ynrHx6Yik67ragOBPfmo6snPLOxbdtqkd9a7wiPQOfRKOD6GS5fCvD7CrUwDjH/ZdnzhyNJ3s1zv
PaTr4UaWCQQQRhCzlZhdV8EJvpUM1WwZiQeZ0qsBsRL6sIZDbOdZTdog8sxku3MtuButTy8BJvQQ
sAsdXCN0LyYu1o+tArlvewoaTmKN5zNC2R/YDvYz71JhPdkSCQKYBUcKVtXvy2pp3ExyocXQXI1r
m5BXQj939tv8MepUhyDDYQcQ49dy1KoTHbytkwcO3SbpirIqsuvaKSreyV2nVNdyIMFzT+TUFkz1
tj8RzQG4HO4pIxzsL6u8RBtAsQES21I4/kQp8uKNg3Ckdn4cNVrsKhxRCXF612Wvber6RIgPwOxC
75zMp9UtVo0BeTkEY95GvE8UmsWqTnc6Bi442i0UBv6BfQXCwsNpLAGxGuTP16nnWvcj4lf4hu43
HPvkLVR5ERqS68GNFIX2rgK6cCe6eQ33YhgOi7x/NAu+/S7u2Z8NQsjOdD/rYFekUXKAVaOutV1E
d4AwX/H5evYeO+oAx2Ze2rYTjxzrIIZQ3XWB0apIdRT61aFIXY0emoqnMGU9FgYGGLyU87yEHyZF
9y6fMJxGLowMQ+lwnl6w7UQ4V4biYPLOfZdi5wAzA/s0G3wMmuodx4sHB8l0m2KqU5CduRtGQ3IQ
26t6tVPgg2fgz6fKWB749lYVWXk8ljHjVi8vO69zXmjLQ23Znj2Hj9bo6a4fikk7UFfKE8casjo9
C3aUOGGqAs4K0/LP6z1Fe2BkThKmb+kVNTmZ5sO7mQSqHpvMGm3P9ybBD//YoziusFmri+zQUC0O
jiE02QyELsnwchwefPwsRCit678J0+pDIA/5XS5jawsgkOuAESCvEusZ1Gv8Pkq+Ba7/ku3jVV7g
ZYOzLSKWkbPDOWsTualPp/OgZaRnvFdQrMbuejat1/o95DKmUxSRPYmTzCAG2JStPrcX3/ZVOel6
sIxzJspczGitkWA1jzBqq518JCWlrDopZ3e1XT1Ed0zUYwd/Zoqa2d4DLMjjAq++tnfiH/Chgeq/
bxOhDK4Smg48DCKvUEltCHXidsUpVaXsIiYzOZmwwDesKoacOmym0HppbXAzeIFQVaRhNbbMn/Eg
JacV8xYjqH0myYJq9JfP7Jr3kixQPbk5MY8L8XbEwrDD5L9u9JDKs5RCbPS6g887lGay8LYgbjgB
SKBQ9MrpLCw3y1Iegh8TkZtBhJvfTTg3CnXoq8GD65LS0PiJ12OhsNgsgfvofZCB9oAGrVy2clN2
XjdAvv4IWtDrJcQmTHasNXBUQJbmv6SB8iO1tOIip2U9SyhhYV5bX+lMsBImTqSjkR5S6dbTFbSW
sF2+qXvtcgExFX8LqQEABZna05TZ4LPyWCmt5lLjxhysXyY30UkDk3Yxz7LrI3K2LSgRJElBV7eg
VEYIDmsF3MmX+E0MpRe/Tt2Q/3wp8589Mnn4tavgmYI8vXLcRqMBthkNybXF4l5xSbQS/I/P20Jl
+IZN5u2B3O0teHlaqvXKwLuGTbLuaVxTqqmUW2SQA+rqvDpRlFxKxdLbfPy/ZIdAM2ClukaAZoVa
ZDYPeXcc2s9XWjxTpvyE6Fs5EfL+VcTQKdzgs4jWxTOUxjfNZmwwVrcEUJakfyv6K7NBfuAx6Rv2
K0vwBhtoiKlROOzSvWuCXxnwcVLNzFiBqCVpz/C42psZSeIpIRBt9VIrlSqW43y86ogRMmtHsp4L
sB2DaBqMo7HR76PLGZaWdc+VuTw6WHUPGY4cWzjuYOS8VzWqlsybpdR4rJ0P2NO54EU6msSZjzVS
u/0q2Dim3NcVIGEMBHW2+nhVxn8eS6FyOG8vIplNGmyyzDfCDkLIMLg5ilog/tnk1Nql/guw4EEQ
8Y7FNLNdyeAitZGmIjCrSV7Xi0nY/b0dqHbGEwLHR/6IIjAAKpWty6HByVXe73UZLZlaq8XP5diP
8mTNd6+LJuJ+1gpL31S537AHlWkwsCPnb5R0VldOe9kGOf7FYnv5fVb/3dZBgdYJf5BgF+ocwvfq
MKUAB47pJmBV1BhpwmTuLFwOQjHk++cvjhvPkwArALtTHihAYwTgXbceXyRX8xhAbz87Cj9/lAW5
inw6gAkjUKMscpU1ybRDZmVuRtFWIqMiV5E+ZiyCG8u0lKCHTb2rxb9b6pEZPUSqn1GKM+RjWKNW
RpR+xrLmw2j+rLESqTaw/ZU60WLT1V32a73gTqdixZpRr+GphWIlLhJ3KWvJRdL2FF2Xhiq9Ji7G
8AF065xHmjkKeub+V4LsZ1viVrHltGnbBFl9O9Bblw3kcpDW3REe86RnC9gyoobKGy/ZcHuEjZMr
H4xwbu5QlzCH6q93jxDo4EStidWG7cjqe9pwLmX3jwC7F/+zx8JYFU3DifWwd9TaB/SAcde+ARc9
hngwgwYjnPAqfRdCoWkWAtJNL4c4AaOWgX7AyGXCzOabqAi5rjtNii1XRcHgyMDeAMMT9gr9id4G
cVh+kXt6cOHN+d1TL05WMyFrEyns60IahNtTVC4V4JDBZ3Ah/wi8WioiKNX2Tfimys2o62oj+czq
CbjoBwX2KX6jEgNviFtP7isWQi6Vzh+f67qxuOpppihiJo4PpdTpw/BqLJ9xamcdxvtoYgqRAHRc
93t5nSverZf03Cjok4s0yN4ePJcOE+h1N78ACVEwMNklf/Jo6jTRuBC7ioeBv3Y6CZdhi4wfEDq4
IHA3Z71j5yc4f79ijw9IYRaLA3HDeO0A5s549oKsVvjoHTyulWfBYgibPn9ojDEh8AMzhxt7txrR
/oXA1P+xbAz8pEGWeWbYeHJuMpvfQcArG0lFNPpRCZH834Ydnw++o1jSMLjUZTQqaVHijfkQQztS
pyFpNE4stRoQW+DpRLWoiW4PSnMozgc2uwcJacPHpNBV7i8d5/EBR9NPPEIMJvrk/thO4/jm5qvS
z9lG/8j1HEo9nEYXuKc2j9jRr3zK5ixGuc4XzjrtvF0hzlhazBMCS8iJK51mzrILZKiWs3+SraEc
H91JWzbjxXIesAZGZRRtg529okRNZSzVvb5kHPdb5zsKxJ58ks2Y8JI1Emp4xvkmiLNRk0IL6YWd
yMr5rl8GX6T5lqxH0mgxgseQcBn8WAwf0jSOETiiXKQLgJF0cX7x+p/Yy6NGprjWg5KdRuE5DnFl
RBTykxDL/csLcW3RhvJ2x0WRNABy9Xrn7t0sMWnNoDJgezQWM6ELmdx0Oz80stMILNg0l2kmdAW3
TxU78wDhzjokhlSiQU/WNir9NKK7QAaATQKJft0VMya/3C3zM6vBAJTXcjOU3O6S90WqMjwVWRIC
CkhJ65eun/PFQ3znEDpQXtC1wdbHqeVM8VMXqGRvB5NodnZ7qg6DGPwCUWklkal5+GzNt6TK7lwy
s+KdZhJFCUYDw0gnxFH5DEJcJ2wlwHTfU84bwuL98/oUn0zhRrA+JuArQDo/OSn4GLJuHVesNox3
ZAgz72HBuIsk64mhIkFVpgFIMZqjdVDcqMBFsDTRF72GWZtPDfNI4Rd6rsCAPmyXL/BbkChCnWcA
6HvQC/qbuOTcOMhFts0hFhCluJ6jqndJxnSLl7D+Tpwb1uK+XpJGHl0feDwqA8KAofH6+9+/dEzb
jAx8wnzxa5miE+9PxgyXH0D3UHs0m9aBQu82cQfoF9besjL9twBEbiiK5FcnDS3UjfzkjYpHz8US
P31WADEVKQtsBcl9BJcswHpOXyt1PNscNDUzEbXuTZWg94NZ7uh8n3OBbg7ut32oudRrA7gyLiU5
VfvK3neBzogkwYk0meH5sjNAz0JyuXd2zrP8DJTKzdg5UH9+8ItJTMTcUEzVDJ+9QUpuA2K9E1Gh
A1pHYtHIDhw/VDSNeqL31fW1lcdPdFDPdEZ++5XvyO/aVigzjmiwJBw53SDhm5Ok+RCpCej14gmH
jAk9tOv01aRPinsU/kSmuyg91mhvTgrJEyaa+pkdIxE62p4DDlgjbAV6Gl4CopyiDO0EHumaN6NU
oPzMCNVD6FDsYRvCnI9RJF9yU//CSRphS7DTFvcsWSvULu6J9+uHI8dtuQGhyqxspN7GDShm36C+
z3wMbz8GTSD+OZomYLV9RYeoyr32z2N+4ihhni1cVDWLFjDiJsHaN6Qmb8NgmyIgfz3DOi1ZJMLw
Jml+tRU7CeBietDE9R9C0mBpAWZLOC0sViDPUPU37KvLjhuym9FACQ11srL6lJCfxSdkMkRl2Ps8
HZtBQ7f0OABHsw/PSaqg+5aB+5nybpLu0kb+vI524v9zEwtWUnl4Bhe+8RuPmNzJt7+YUm4yooVg
VSX+Fe2An90+KMVPwJ7ajNaZpaAOBDn4O0NqGbOIBYLgGAq9tqNWILG+GXSvpGB2VjwNJBSKfzPj
Pf0MovBq19j3AqOgKFJm1RW+CigufjIXeO8ziV9TWQaEZqHp0/PH5x2EWi2w/dX5dK/3u1lFhQWW
vMNkcWcq51ILtPhpuECbTZn4Xku7e7SJV/HEKZNz7NstLEK7mZQwozt9W6+yma3pqtcKghJQX60Q
fsPOYhf66tkTc/+MUkRabos/EtcUWNdmYKIABgrRScKorLtaHalYX5fZqo5T7U8hyr/QkDdp4w1J
o3HSuBOlsYCpkT6eOU5l8xskopt4cNkrmqC4qML3B0vpuqZJ6xtPdqsnv4rQSNAVk+s407N0MhLa
sb16a2G7LOvueXRVJazF66TIoc0U1oIxJHY1ydC27Tlk5MgEy2zYk4NCvVlRdzuSZSg7SpphggwL
BXBwQmbyPxPMAitdFN7yglPGaSdyL/K5Ta60zsKdoCm/1dZ2BAY42np40maaFVAyPML4dlGixl7B
weWHCWYepFoteZtvSS2LT+X+VHGkcBvzyu6LAiMyz1eouUSNhnVHkQ4Hfj9m/ZYtJQ0Zf+P7J+wk
y82lB/K+QOIynKrz14UfOSJhDyaS0efgBSvlMsjR0KJtvDOYF+/t9Pb8Su0uYtgb5ppOZuwN3uog
PUOoTPWPUzINrKX+CD5qoG0g/o+Z4GP+hhYWFIOE+P6ZNowI6Mn9pCiYvbIQVikk0DauvbKJcE3i
ADG70ZA2B0sClzyxyi8nJA7HhqzZsCI0KGGl4dac/FPB/f9Npxw2HdOfuhttYzgS8//FYjcfhYdI
Jq6ikfAcWgBIGqthIwjTYRI4Dcz6jFyfMNF/0dfM3r9dS/IR73bdq90POiiv+MHmbs6p7RoszXlv
04YQud7VJAcZKEY+7Y50pxtCEnYIHLeTsTfbu1FYhDyjIkJWO/QXE19TZVwoZ1rxJEDRZO/8sXT0
tazmGrkF+3OgaWkBbrqeb6mqK0Mgf8DvPnPZmRjKNO6Iyv6sRqZmDGbV8kCmcIh8SFHGQxGdVg5d
7BP/mC72C+7vV7/s6XnB8m/Xy8JnKyuCJQ/Bvm9Ppt0BobaIvr99lNjW0mqIyzBKMTAB9xaNPM3h
QJEgMjmLgB3FOAUFPUOvLxi47F+wdjzW/q+b7SRXtQ8SGC5253vNBo7jjuD4SeWXm16MG+01y8ZU
tKGW6fpCxVGAkBoytzQag1pFqnEoWTFzqRB942D9IWBgHpHYY6grjF7HY0lANcPj9DQNrmeDMfvc
pLsdIRexG5RzwzBxP/YFsLA79zDS0IAQIsqk+islr8ouv2WIlukqp89hDBjau2ebeHMtfbpQtE6k
jyHs50t+pJhcaCAhWCHHReQbVuBYaR1Tn8nvYfP2n5m6g/ZCEQ+ge8rEXyWvhOy6srMZFBa/rzJ5
pKNF4cUUMo3OPkkgdZCj868A71cP5DAq9DSb3+FwLSESY81LBiEzB6lhMlceSGMOwKNl7uLVOAUs
0aYmsvKIp9x1g2KX8LokEb3pllQ6AkXpOWBY/mA8n6Ikd9EnRSzPUjRJXl1kWYIdtVmoOkpxpbw9
xdHzTqfgESPe6W4Z/9WbLMiJbMKlGywRAky7u+548jMo4gH2zYbhYZH0GsXqCUzEr+PMe0nM2Ooi
t6wXL/oyHxs+UxOT13bBVwgWoYSKhGziEyt5QZbVwal0HXcgpa4eJolzUZ17+Fzq1pK1rgr15tBG
IM5B/QBCOutNZxg+L0G9zQq4stbQiZkCinIoTZq5xfZvY9DJQoB+HmAp5hLGrYcPn+o8GX0P71TX
/Jb36kL+xekRhQtHikbEPa++5LlUkTgIk33W+8At/X0SNlcWCeEQLVG7UtBL1FC9OMiVsYooZqlX
Focapo8kxlbEo7LtjBa1RqXUC08untyZ3n78C17fKRKsIFqgIKiwgponrzxLvIWPaUlBFdT7YgPj
FZwmiQSPn26LZKJb+soAk+sBDTbULJzgOo1re+qj1UaDQOudp1S/vBtMubASt1jsIckwgZp6y7A2
QpIB8HwmATaIby9+1YbE9YDauIQJYtmSSbEnHrzp4gkmGVcnARxlZvQqMNSUb51NAy/cExguACyU
JRH8qwvD8yBwS0XgjRbBStryNw0l9CYRXhU2qcFQRBgTCoPPiw7dB2JUCBGiEvLTHbEhn9mMfBl8
546hRfSnkmOvGz8hXeQ7wo8PKDoQHJsecPViKOTOAxueu4Tb+F7dUqGjcG3/xJ5JrJxrvztbzWFd
JI04tQaFjT++YB/zjOTPNYPZ37boNGrFWEae/+G9OaD7/okqSvkW4zQOHELiTIGhtCLBiGD0NAwS
BQm48PxltTijLLSlX8o1l4sN00fg+8UXQlS3vrkx8XnOjF8/TfexwGsxcxtUB0Mu70KoZM9tvbpw
Q7Mo7tZuXUSxcbVZ8Nge17VetRJ2jh0Yr8am7/cZAea3k5Y2zcV7b2FIcNl50NAF6LXAyfnzqsH9
FAyVH7ZRFg1pahxqErQKnumWXSXd82d5AzBMhQ+PM7MBAAxiHr8qdeOyLfklmgPgq5gkdUIpu19G
8M5mPTBPDYrb34pzymWpcGbhdWUaVdXwZh1Lu6/tQ9gMJd9t5LXXLnLQd+m6Jv5bL7Ex2vGom2il
iTlka/nHCGt15APhmgHgkA3PW6dnF2gvxg7n1JjmisbaURBOQTHAKho5278QupvnPOB1TbglzgN/
B7+kjIMN/gXk8InstvnksikHTFAYsST3SHRip0CNwhW6rRAl1xh55dwcw1kpmSIjuSk7AJKBSs/8
F3c0DobWxD+937gLLqgXo6bEMz2j53nbrlJEsYMVaNT2SG0MWD8Y8HOzxQYhBe2AJBYoV7JtlFh/
oRiUXBZB3dVDKwRT5mzVtJrMYtJIEf8tWVXrbAeZ1GRaRe+0KY/a6CwbVgJjhPpiizQYeaSGOpPI
vGa7AUNs1IIskDpmhc5XuInW9e7aD8J4yewCvS3weNyX53SUSEj3TzIhmcpDwpfluiH3qQtjexMR
g0XdqSXHmfppp3cWK/lxJ353Qlmcft6kBJXxAyWUVBrHaaMNw5NEJlbMP0ip507AlR6ToWMj1j7C
Xh1p5+0NLcgmTUPVVlo2ef4lyPCpPHNin5FpXzi0ILBEUFJIGPQV41s88QR4e+7cGtcgh16LbIZU
sKCV2EpllsLVXceqmSozfT3TGLvVNp7YX8BneSMrF28pwQ1w7DdcEc73yLWdEawUCV53ZaV9xBw3
XpHpnI5ihGhcxggUzizkl5saZrvgp0eMpnGjMKHK+K3IN4yzoRBycVl2pDIXGiHmVycqnH/moDOs
y29CyNHcMZcnGjCcM+xz5kXQTv2gpeFh2EqCCYQs5ScUQ8OWW96gdZQs1AxsESxKTqjYur8HPJ9B
B4maFQfF33bk/joWWiXOmmK3k7wW1pcWLOcFZaGQjfGgSJ9+tsDGEfBpa6WUKmPMoHB7stCwwOyy
fXzkJHXUMZBGtzW9mgDtzTwtFB6IKNaqL/gfiQrQBYJTzdGnT5By+N5s9b5rZebg+4JxUW2Xdl8A
oNz3y0ASjfkXIkS3I8KoPm+8sOpC4al1S2eavALmB4K2EIdiyYpgubHbW07Wn2XZ1WWRpTtdWbEl
zSzHSaoPfIC+uFj2IgWnMxQS5faC1YchzhEsAkZUOCdbIPFVAhQa5vq5e2xmmlof0FBrzKxJn6+k
sALjvzZfg1wMox4icVX54Z7M72xLyNZbwza+CcD1299sggydeGlOmP6U+8u7pK2zvTTRwaIMV4sT
73ujTHEh9XPU3ZfntOpPC6NoOQIXvLpzjsj03O9rzRrmFMWvylCSlWqtmOnuUaR5lgb85GGF/l0Y
Kvssyfv6+w1KgjyDQ3mFFQXR7Ult+jGDMZ+Z2VvstYBigiFeazHSY2oxyAOmJRzl/4pXMA+pM1TT
1imui2fSgPqphqY6VEnys9pDhqko37rm2uXicoaCtxHY3S7ortfCp5+jciefIiExdeqn3Acy/vUv
e2ppI7/EnifhKwhc+YPIlaPJfQxUbjE2/BjFjKYucS9qe1xlSkLmRVU36xx7VxEpEqu6sX8QdEIK
PhhIYhPHh02wZO9eRnaFyN3YrQ5u/DvQaebI9Kta0YZJEB/r0wUq8giB1LLxR1IOJouIuCzrQTcq
DuMJdVAomzejyB45Njc+DnKNqD6k9ZtsPLSeTPSuGJVGzFITa4mW2G7YYDsVc8JPyoCz36PQK7EF
isAsoq91BpeZ1R66vQVxjuUDitrRRXirgncZ2zKRpjIODJ7RL22jXo1AYD4ztwL6g0YVx24ZhHdW
18eiV/iDSRZkvi6oxCP6X5SytGQNrDs5pttWEtiVfEFfBOsRGjR8zVsJcZD8HcFmtum87yn2tJLw
n3SpH4ui3eoxDkgWc0JYIqB5m9tYa3k8IeaBJ0f2o8xMpqRWUx1an+g5t+qsoL4opEVBr9+h0pP/
ITlno2Z54muTKzIS+q5GiwQoU0SZVpA+NcyndpcSGNYJJ8XEh/ur7tXA/LsXPfPQY16R5frydKwe
VlRFB3P1GaPa1RPueC2h/fw5ni5mUfwHW02avSMKS5ymDQVU/FFKDtyeyJMYjBVzH0uUTLFdpPz9
V1qlyrWNJS2gm/pgLqpjQq68zeKzDHLECs5cXVCzME6j50oU9395F0lfuvb6u4pB6g5IvmwrQ0PL
xuc153AWK3r41wedPTpxgrC6uuTk/biKyHzToEGasPO5LSbMXNS/icmLrHhgOSzPwu1uHPSNWea4
yrLLeH/U6G6r/Kysu8sEp4nUsVFQ96PY+P7iG+Y2x5WnmCGZCVv+F6oM+Vn6KFvMJ9YIEufZi5IV
lNdPWZBRYujqTCK+ZiGVTZ3cMoAsFoxhlmUN34t9RvWXAy701T4iZPk1t3uRh6ND1zXnYUNvHtrD
odvaQyPHd8nbhCcEW7DLlydXwLWCJsuuogP8pCapo+flPCdoRpQRJGOQrweLurCe+3UrkmZj1sn7
Ot/zS+9s5XG7BAJ2L7C957B0RaZ8f1XmK9NI3gWPM9S3OXqMuhcESJ/cuEbgDG/s2RMv03kYmm4d
1e+anVFMcs1ur0AkcgIBzZxzm99tpaw24QfwWBCbNTeF2/0dt0o/QvEpNs8e7ETn8ATD/lUrLKKp
abHsOMhyANWmZd4v2VEcp+KIRXcXBqqNfWjuKQuL2nf+DwJQLVEAo7r/rqDSZUC+nxidw0zRfCAr
nvKMCFHXlfJ0pyQ4UFT2AiMRDAn5C08/BXiiQwnERGzPK/mhl8Ga0/oYiDA0i1n0LHznKL0CceOm
NfEfqSKAXcMfj16LjyE/3NCIolZhs7W1pPTyl5WTSVLUlg0t32Gl/ACSFu81C+4DZ8bBmNYJR8/m
t8c/Td58ittFe90NLZ2hYManh69g1Jh2J3nFwfWa/+PcHVMcV++8VzBnZvd++T4bJCr2KCtU4H+N
5cgOytZ0OcIVuzuGSShLvvX4VTnFFCjijhg0ycoJkX8G3BIh9hxX7LGRxmpgvGI9QMMDYup/z3T5
H5UWKyPBqB/NBl8IAfOY5+lUnc6YP3pClfRzDO/ulrNwfKU+f0P6Nitpm51bhdUEl75p0BdhgQCL
KU0KFo/VkllrqduM8Bz07g1K7flpBqlnWySWuB8ALBQiBOslxik3IGSrZTbYfs6ByjoctP+L9btv
Kr5pxvBDMRCvFLZjxHmPest8VRXhBIHjnkpJ6B4Exo8ZFPJb1ozJh64BFexrlSdiaHgMagOkr8lc
q1YduZazY5+hrFok87jzvqoKKO7Bkm0VVLZGh/AmHmQa4rFxhwC6gJIZxHcvlGln2L8e5TRXF9Ao
TZNiy8I7jqvP0JLp3PVPy8gzcs22R22xBimOnqv+3Jq2qC4XChr8ZOm/7uuCEpevOy+TK3UaahYB
7tJYUWMwJlLmH7+p7RAd93Y7zSdbit/MCa/Y+NohcjtKeqMVvdFwfYptDeXqP1oPdnXDsvLnWcnX
cYNLgmBOXIyO064YC9E62/UiePFBKLTLevj/D7JxSBe27m3qDktmVCz06B9iuBjEzgxZZO8kT0YB
2y5r/SzH8lte6rIqIXVBaxUhu+fs9FwZ8hE+alh6vYg+c8NMwM5IG32wvLK1B1fCmoXBaDrzntwd
rv8Ri0A8SDP+1yuQ71NI7oOIqBqKPhubIMITRuEn0ZZg3/Y5k9johVt5fCskOAET4+/4qouQVQWv
Cw8xBKRKGiKkXLh5j+R8ckLie6TxzEqqM6DvsrtY8JHrDrt9hs9+zSlOijceJRHegOVdTdfXzN0l
rSvVv3nb3BnFtbKMRhe2757V80hLvCbLX/cr418R3OgJXrVvPH297WpwhH4/4rn1R9pogFa6bYWB
V4PD3BnSdW1cziUmciDTJzqnmS2kK9N5l6G/hEwmYvNGVt4gcv8IjPDNH1mWwy3+5jKdAN6FZbhE
COak6mzQJWUlD4tZf60hidW6Ic5Uxc5kjVsfKO8XdKPW++z6u/qDSaXyBuP806cR3p8zt074Crdk
rTJru7xsRa6OBI+nCNlhGF0BuVUmK/Z5vnroCMoY6JuXmPtLCMQCAyEUYO+NIEqQwCxcH4mmdqNj
4I7bYLmac7sH3XgNI63Tdm8VSn4JPsjz8POc1kL2IxQ3wmIHV9Y2hePIh4s8b5hWfuk5yJKTjre5
GLldlOkyngq3OLcnaFl7IS0l0rcmbQPiJKK3t8L7mtUsCZX7B7dXkVbK4G5ZyEe9qRytYvchY/Ul
mnTh/q94xfWcvoPi49Sl1NPitmHXCU8P3M4NAfh3PLuYsUfwdTnjOccDD+q5Vd+pPaSLgPOun+zw
W6nJKDeNIQudWPaBjhAqx3G1rnTJXMpTMKf+9dmxgntZp2L6s/c5Jb0Gm67/0jvdHOFIF3/PehsJ
+mqcmy6zU0wZA4EANaeU5lu++vHc/k9tY6rIDs2BDrTnUv6uRpuavy3qYN6CBtn2JfePdDwqri6i
0o+2SDkBWSyO2YtXI73HOaA874dJ54bz4BHp+L7WDTi5nVb0pG6LokuYw50PDTDmxYG+PwbBND1M
LqjFrT6OqXLjbdf4MVmCYusABWhTSkTRf9xUCpTlUDkuHEWgPQ8bOPh6SDGqitty0l5VwEyllZ/F
9yXnWAhZPIeHlMpM64E6erDTZZqrnC+5HFmdPizWDdvYQ70MUn99Pz4EWKZ+Dd3GEw0FPJAymE2B
5qYw0xcRQvOI0XWqGzPhN1bRJoFP+MQDjeHvJ0QEccGNcQlFZIxZrL7fk58TPOxxd/701HJjek0e
R3ZfxA5ovuT5W6fv1odPzF5aVlFbwuIiYCW84OLcxs+UzZJHXBMNTcz7woOQGJFmlNeLLAOL/4DE
+xvGeTdniMu/9+E3yGucV2cR20hHlQ9bm63ZNBurN5vYjWFkMEM+tAtUtUWyUvqLyR9v7nJG/koI
8AeZ+C7TYcIRiuLBthCW9AuWpWRGVnkwCWjRXfTvdx9QvdGPML5xfOlEPKKqoZZa7D8Z5fXqCbE8
XRyMSzzgLY4hS9ocUwR+Nvno9PJNYMrJ90DybIU2qMrohY4ee3DSEk+/y9jWN+1Qpj8mF7Fs4dwv
K02nUOuYWyAuowf5skhLAi/nnLyuLH43CS7oNxM0wMn/7GmZpNYvI+SdnoOEL/5zhRhr7XZHN7wq
3VAmsyI=
`protect end_protected
