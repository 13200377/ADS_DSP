-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
sT1D8C/wBUKL7cDu4jMgUAWpfyvsAQWvuk/nmwuNw0qD2SJ2Gg65zvDUMBk8SlIs8sSceDG//VfC
myAkvdfNeQjrg5enp1k6Ugo7qx3cnSHLHHhhXN+bAPcNkgGyxiSxYEtKI5UqybV1+3gQePQY0umT
FdlSXyJclTvzWDTeddzAqzIUSNybiBd/R4vTeFlr2VuaT4wojEapYICAP/OIxA8V38CChgP/Vd46
G5NmRX0YeIBQNFvQbT6tcsAcQI5yHtfCXLoQrOFxqJawOou+w11/sjPHVSo9Zte515uAUdxiL7xN
mKvWrUnPn0ljmvNvzzY3Lz6Thd84OmPdjktbeg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114272)
`protect data_block
M8cmXX36fSvlST2h0vvlqvwz12deWPqrEkeu+VIl9k9Po4fccR6elqw6fnUC5X9x9ix6atstfLPv
8Ot8mLJzFruJBim6YKy//qXfG5vPk/Oey8wnWUML4tQ6yF7s+63K0rSxbpdasFFzzB8qgvVtd9oW
eggLUaABHNqPalHOTVhnYTQByrAjmqHpOaaP0biImUARB8OYj7tHu3GUN47JlwsPmsgfGFu8FdjT
B/B5zbNVODE1uSaSl5YL8AXjPtRASCGncNSJYefc44lHjvel5WBJbWkegXo7ddKgeJBCt2Q/WvPD
DSXyv0N2548nt4rY8ZkzrKQnFqgXUamIkBc9fZXYyc5NKlU4sNgZJQJKVCQm0layaNIUlPx9jU09
ThSQxCT/3BqP4ovVz+Y6G35UNlAuJeMI4b4tugvQLTJqNWVw3fO31Lk7+inYG2HHRZ3Nbj3Up30W
sWuAFb7Cp5hP6w2b8wIIyaZcJRWrVkvw2uwkilJbDn+AAIHBB1s5zZOgPXvtpP3ebqa29uJZLHUN
JqcX/4jhCT3c2sp2ieEwEyHOzc4CfYo9iFyoKRHoTLOCEKU6pUHSbw/oh1j8yCnKwQrEUi0F471b
DBm38HwwT9lzasYHp3uLbYdFFacLTY99vMuzuONZ4oY/ixuiSwaHoWDZ7FJj1NVCGWtVE2PSYgEO
fI7vg4sSf/uXsk7swGRltcnHU2hhpfAVCRnvUV/c+BAq/TXAgF9e1BMUjQbXoP9As9XI4YrNvTSq
/yMsRI7TLNYv9qHpwjnTCKswdhsKSOBIhn7fTcgQcgL5KSn+LiAjs1d1sEwJ0FCnQuZFIbYJFDxr
LTuLcP8B/enknDv7ZGLy/51dWaW7tGuiYFlUwMJ7JmpXyOhO18zl+7teA/K5FXqPvwCCYNV1z//K
u7tejGlrgAFyTp7HnsITDnSIa7ntEWXwlpb7dtz7ymyf/y8ZuNXfnh7fFuDP+tTiCUxJ27yAY/Xt
vbxYD2QtpFB/RHfRAJb/0gwvUAuzX/QMjv5yeTf9fa5A5LCkiL1gIUbogvrNswif+tsCQ+E2m9mV
Jxw9fg3w1Lw1GWxoqhSuT1Jkfy//DemnA7x6wUcp0TQxXrNzL3jeqGfEQiYF5AnL8FDf/ED4YerV
ZpRlUcsVDR0HPqz9b2heFhJfLgI/U9kLAPn4Qeb5K44XX4hbMZTDfcVYt2mdsQu/VayFFF0oX3OC
m6BSGJL2/uwQay8zsBGDur5n3njfsBmZ1whu4RNB51rPvK17VlfdgwEiwBIldiccq8/wjwyeAWZv
KT5aXby0dcKE3L0YhUb7VYaFQPS8RvtoD9TyfZA7fT5xB9U4575MYFY2tark1BftOAxuIU/OvHFS
dzqUEnQyyIFfcUXelQ1SsVSefElWvHGvxMEc9MPsjtg4sUZcpSoAjg2/wuOKLZ62+h8pHyjW2bed
XaCfDWvG9/YGhYOgAEGvH4AjFK7rrJhCOg+OohIh/TdkJHu2hfQxXMe9hbgbqemXgkQR18k09Wim
PZcr+B33oC1U8M+sNChcRfbtabMjSdJZuJjAB2KGSfraF/19E78Thfw8sW/BJgKofzkOZ3YD1KnM
TkBv1oxXQuJLPEx6OY6EZyo40v1StTtTTnKVeAnNbu3DT1i09CVNFg9oVxScuNoJlwgUWwIs8F7g
wEnEzGolu40+OH5x2ZA3PZ3oSmBeWeiGeTgxrHDqTAM3uYHud7SfV+GLzg2LTskeaWmCLl67C1vO
32Pgq1uhHZTHbiSk1TiW/eN41Y/8yKz1x44gSz2fBBQKQ8jhPwDO+s0I7GMNcOluXEjU2pex31Gy
/zJ0X5BSrP8iV199wf0ouIJ3795kNJB+j7CB4rJejGnDoq/v1xWbRDC1mBWMap/q0tAZ1co8FAHn
qQXJegxp06pAi88Admjn6BE2NA7wa5gB57B61rWvQ9M6U4/xlL1nmPkvWCl6T24TJA+fJjDLpGV4
tQ96nengxxDH2F3snedpk10Z+7WOKcgz2peGIF0dNE4S8nLtDrIIZpAhtoswTRGL421Y/w1jHKSd
CGLLeXlz+uIOU7XiZhsJ9jCvS0Wg6+q8iHapWRfXiJYSS9dbgeg7DTYQkQ+7XBkkReuUKXl/KqAa
zKXSiDDpVJQtZjo3FnLdEuixBNFLwjEme3A/xm61q4zAPuACYyxFc6hJ+dC/8hOVKmOLsaC/lzDY
gYAC4nYqP46w+ALGi4hlMb32lD8lCyiUR/9uu3/c7horYNmUiquqp6fEwKwWp5h7+ipQc8RYoCv0
qm/UF9vDXZqRmJ9hODJmGU2GYEYGnNe8LazjxRXXkEjmcOIbZVWNg2Punp7LQn1ZYuKPX8nqaZO9
hPuEuSxuhgmWRx3R1n7cchthaBR+4HQ0jergNADzPXSs+mgm47+vcMW3HH0HVRB6tt58PALdSQ+6
upyVWE4ERx9vsZ2nlan6TrwD+8etjJJPjOw6A5y7uJo1FurcNI6K9IvFQO7o53Bl2OkTWpBCPpw7
OPxFgtZvcveACp0BWqNbwQCVVD+y/fOAGY42nkUpZm3engwCCr5us3gHyoq5eTyjbFu0DKjU73/n
HtD0R9mNPDDE7ape3yOd2H1Pu1lsmlIqtZc/isx9DUsThL4gq4PR7nfl4oj0V5M+xtYjMAgF1I/S
9GVSxxtqWUJKB3ORHiKcoyFZDGGi8cUWykV8393cKoh2UxzCZpwsovs16XBxZpIeSHC/JZWtIWzF
xWFC0kRilvKi2UcGcwyb+wOyK9O05fQR3MOaZN2Hiq2QoVn837Ok0zOvnIFbogg67kB5CVGkBK1k
YriBCucMlunJr1PSoStEzjXxHT1vER/v2ZnkkIGZvPeqg0RX/1VxtOW6k/9+eNsZUJ4TFAPnA4ZW
SxYX7UQNkNWs8D9zeXOZ/31J/K8NPwkddqf+ND6re9qWuHUcw+6O7Y7oceHWE+GR7InH35z9sMa4
21pKpkPlSS3619QARj/LsHPSotqfSNRxIP317ON+dY/WxLf/2PKnpHFgahTrG/R8yQlFGgfz9yO8
wKAEhy8PHyiYqXynCLp0sZ0E61ZcIrgSVTtYxHmvfNDJ51GllkQaY4HVFeku0i2Kao2maSA8kb6k
Z4FqoqTGsXQfbRvB+uZAwoehAE10RcRXa/EbnXa1hJ76cdyk07ky8X+yiaSQPmvL0kGHi40JRCT1
dvyJK+C+WC7ARZWSLOIsqW49dt0sfl1uJXup2DOftXhrJFZJah9OjgRpmzSK5RMbw1N7hlk1DMzD
2VTiWv8XVL9HQRrelPgG4CkjhEY8zmhGu6M2X3OOTMOw0y9kF7al0/QyzjBOq2oacfyjW5u0FQG9
Tiy25/ALIFlFZNlNG+9/+Em12ihjLIEqVv4dOuffH5rdJcOHLmSB8u0mmMbzDMjlGZNH/2y64hTF
B0vk+EbI1KKuXwf4rRVyQcwbcZvq0oLDy/41GeJsy/OPyP7a6PM7myaZdDKC+W4xFQnSh9ezOcw4
WQwWAePAKCU+Hv52JMb1QV7nJZmXGawzIV0yb143D2Q/p57FZ/Yi/8mv9vgdWnkP+i9mGS91KH6U
MyQD4J0Ln8Iont1z9cYe2P8hg38wUZhgJgmVKlxO7J/YJI0z5s9ksYzgWqJILkzeV2deST3kLCK8
90io9ReJDEIPEMFRfysPnNDx/6/pCFv7uSbDi6FYuHyKGiXmdOCaz2xeHZ4yvDvZqWm82R0EvOkY
HaAT2BGUG1r78G+qpEGQAyLoKpk8Ah1Lg2U/x+tRQ0R3jz+AMONhR1zqgbCmrOPrHJ66Ok6oLg6X
OeZRIMsEVSvTrElXL6mW5NrEKkF/y5KjhzmM7i7n2oleGG2xovTkq+O1N5WlN0gvw6Mg1KbyFZU6
QE0fxP6xNDk6ZXvRSplauNk4NvU+1EYaBKnhi3GXbn4OQ6kCGW3L12BRJl6dFQMVuGs0Amcg6UOy
T+vN8DAjqVRxHcnBPzdWQprGlJIcuzHgWiqrsVekHPIa4BkTAFPmCUjmSBJt9zHPHy5jRBWuiYy5
wGsCPSEeZ8UBCQFWsbw1X0T2gi4prwqNYmGNEY/TfT3A0oaYVGJftZNQR3PbhJ4pnMeCJGdJlcJx
oFJMm9LZ5O/Hj1cknC/wHsKdsIGiFa1Mf3zdRV4hfcleD2NXSSLSe6w/R4YeaE1Rdt9Gq4QFNkEc
Rrmz1867SIRAnMCfN50SPSdL9CNnqXZR1al86UNuUv3ngGONRNFDsTod+neb4e+vNjnhTZzw7ux8
4Wfb8ktaGkGAy43b2Tk8rdWkaysi8azVGX39G92bhfKWSNuAh5PVSy5OvimQ+psoaA5BQyob69V8
/NUhsWY4hTv35aF8cibYFVCYLxD+ew+5hgYn6bP4A+yc+J9eXIpdkE/uDc44lFdAT5YR7cqfky1n
RNPV2rdKtErMFzojTQ8Ig65v1jj/HGfkch2PKcCejBySDi7j7gqI7/NCRjviFcKvh2C38xfo7vgk
rWcaTvJnS8gsW71UDLwJI9RqA+xwvab9VjUw78hRwmwxnMXhDRol7sbGYkSYEWhtTnpVStSAz59g
X4hyQ2zu1MYrkFFiAJ8vBsWG2KnwXVwtkz32EE7drOmxmudTR0ejCFn5mPrgAslKO+HbpVbY3P9a
fFoU+QUxIfN779HRXhhQiO1KRonUBkfWeyF5h0QAPBtvEADeVVPEJYIw/xU+XRaMGNY+DasYFW1q
zzOvksOw/HbFuBrzZLCMeGnEG+7OdbljRGqrxEBxAA0271o7bBsoLr0YSzo5s+3ztw8CHEbNiAiU
zJzBCz3+yBizsLSramfQE+qOTuJAWZfBFMiNB/iJdDyrq9761egvdk4JabucNngwc0rXkIIxrRiB
ShaQtKtM3NKKCduXmJebjE2z8tNk2CQnV9BeKARJ11qu+4lHhl/Pq7ZDSm+hQNcOAKFsPPBboeF0
wKTbdNTM6nC++SNwAxAY3BdGrd5+uec/dTndVKJHHIKZ5XykBqGY5/v7U+xGZw6uxwXgH9DLuevn
0RQGyxHvarghLjc5Q/MeIkyXZ2Pykp74wKodgc6I5L2o3b2eEijZpopgMfIixfX6khWmUmqeNDe8
l7VrbAUC7qn7kbOj2bYZ6qrL6GMAMfPGfs+zbDUqzANGIQhy6Zp2oZoT8U7YWFLYxGLgf6JJbNU3
HnC0mdCMYSutYAELuL5WXQqy3ry35EW0g74S+LGEfoLwG2d2ijScNdFjnwAEhWUHbL0Mo7XOLGAL
5jBibLRNByJJ0eG5/ehBv+9tmJctXgaCOTNBGtD3nilAx25Y0UJbswUf/vMv1W+H9lSBridr32Ol
4R8fT0djSEPYu5DZzQdrns/kAj1mYtvE1o8pFp9ncExRgCukN4CIAKnJrJhl34r/x0n2JEhGf/7N
GWsMFvYVvRIj1K/Vssv8UJBYD7p9H+pBUoK5JKS83pP3GqzhijUkU1zFLL7c+Ea3UnJg6WHdop0j
rePxPlzwlgdpC+HSWmdUp6de8nkC6C+DCO1bSG5nX3m6CNnqE90qnWVIiiiBTrIFlKOrKNeKPcaT
l0kx2A60lp7x9v3HtM2wFsVfcnezSwqsu0/e7y0Oxg3ztq/CdH71bNeGAYbIGUhcv2eb8p792A9x
ojTckdT2YeIhq4xhu8QKq+VygTPe+iWrCROyrRYKw4vGMIiUucgdHfUzDIa/lhGvsd4BZdhaAkEi
xuIUAYnOqKCAX2oPCgThWpSTHQ5C1nzIPVexUl849R9JJx/daXphz2PijdZ+zLgPM9HWkFDVAj6N
AoIwIR1cgu4UIzQeWwYcvMyCmC1WrN5X8FNh3pnPFLlEPqPn3ukY/g7EpvF6CXViOznXkpfbci8r
rzS+myUsvxJ+JkBbRKuGofwDcJngV/V85DCl/0UVkLXVmMa/8m2mso8h1qVma3Ij74+fVqGIzBNM
XoEIPH0EeBcQ63nW5jKJugp68KmVK7tAA7rMffycKyypXIAHatJ/GzP3ervSPkT80kEtCMAPE3H4
63LFU4URXCrxGFigsmxUeTQ2BLkS0CJadiex2v9vb7yjTcLm7pESOhc1dDyYQoiFukMR9b992HE/
yUMvwh16ubKfx8b88kTkzLvtDsxZUOzTjIyj/u1zRV10aah4s4KBJOerjV/l/TpggL/QOrEnmy6t
3az80Ch+/MpnLRBjqwYfBfMLS8s72xgZSnPdmahKxwiWtl3E25JmXQNhymqKdI96KMQlUjMs68rF
I1FLtyKJFSeAaGvE78QT7oUko295JR8OzxwRJnuixOIEdnNXRPHLYya0yugcyL0Ag2fXi6DgSHm1
T0T9vLyPEKY6hZ0Fq76yGt99sgxKYVGmZsmTpvTBOcDUdH6OOzfrlM0mYS3zDVN5xmnngOeUBiHG
HMFyOzBVtYDPVcEradpLKC9Led/lh9nE4Y3ufGHYIiCOln/0a6I5f/6488GDA0jABpoUqk08Kgnh
S7ZvuDjtTOzfhxOtq+pNUphumDh2Ol4t6A1y1S4Labm8te7PH3WM7K40VXb2f/ZyrVakrgAWPcZl
UgeIQRRtl+KegwDSRUtn20Ys5IPbT+eLaVNrwk5NYHUWaenLDtQmfKK0xeMHPF643guPcvpxEl9E
82221i3gOkfXFuCzSA752sxWbkb1V9miOJEOUZXInU7zB5B7VS3erS0WG2sOLoMsycAbqNvwWboP
mAWZTiiHgkBSnLUafBniEkq/vv48izpLyx0hiVrkTdPoasfasWzeWhaqVkbhoNgy8RICQKvpnqpV
jJQBO/k84cCK3exzy3BR4OH5izDXx+CrBq7GfFZa61fOB6EWCiIpvlFj7LB7KuCjimRzjNZCB8ux
FOzdJyT2zLbcva7S3potiEr1XW6NKzvbnZBZWNyQE8HoF5kN6pBsykH/m+U3L1yR5ZsYT0c5GZtb
rTcveu66VvYDYFAxEJ47LJmjIF9n79Idby7DTuQIhuKAwo4K2Yy1vXPq4VCHY/lSprDYfWyhDS05
99IhidmACDIdCtUZKqTYHxoiKsiFqRVgIIUN0y0vMFtHYnM+CgI41+0ezDi/M4YvIGbsc43ad7mY
k56HGA8VubiSu0ewbQy0QpGP7a/sLxOmXOYOKvZA3JEVgNqnR57RCRYcxUQNQ6k73pwtHCyl8XL9
ooz5FEc829i9jX56bA4Fd6EocuZ3sDZnzvanLrnF7EamF4nAAuqIQAJv1sVdheTVTx1qeSaalYpd
Hf4mRjPku8Umclg9aDQJL3NtiWB2H6z/Rqc58Awa/cBlDwRfeV1CCoK8iB3fNFjPy18SN4kmQdXb
iC9BBUlEsQJ9CB0Vn0zQ7RifDMovT8SLjouQSZDCuDNnpgilLrXC1w88Z9X3C/MM6PVKZebH+YbF
SIDVkPEuA9pfUwNNwSppmAmO4S1p1f7mvJwuK0s0C8mE2x+c0JXbEA3qitfg2D9N96oHhOlT7lxF
/oSzLKWc49qhIdnS47znsM2KVz+KWoMx+tCpYMXJwpG1XjfKs7tyLGXma0llmuK6WLbyQ2U65ahF
Ag0MNo8Wf09/K+bCSeldRYWLFTAB/pGYr7RSvGsg3mlY7qi6rDhZWwUTqNMeCTtW2GGOU7284HKq
M5eUIPS/vSDCiVrtjLlFua+4bU/m0KSGc0rk8Ga5PNDDfvSAMKmz78tiGxJRHb9/upKjx71UlmcB
zuihWAIPCUILT7beTssgH28KCfFsW4Zfa/CybKK9YU0oDJGHAeEgMJ+qSoeEgo3O2VAvWZSdDiDh
VxIQ9V4zjKdz8RBQVNXc4ghA2lda2i8iyWtIqyHpfbtzXPL/b9FhDlptQ2wINRldszt3VlCTY/cg
DDASyOvZiOSE7wA1A+zS7ruSsfxBFpFya9VgluWmK0UWMpXxp/Qkc5g9Q96gd7raFrZX0LGJ/gEe
5uV1go38kuW9/LAcq4IqmjUp213PPJ6pnobFt9i4B4ZUt8/5bhCkosipVgFThfe139XBlICfHYEw
B4yDIWqKXOl7pEmtm5yF5kaUqxGf+uEzl6vrLkESZrgGyzAJ34W4vSS0/bXbFIQ2wOxYc0p9JZAb
ckkaoUc+nYA0Oyx0j9FQpQD7Lp6rpFkO4rUZsasGhkCcE1vjUevq8DttuLgDoNXUzPm15ZgVF99S
hos4kWMEYNAhaXmyrEz6BYZl7Wjza1x7NrjiOo8mVTayeyCgaYC/cPlTIQ3oE+wLFKVsy84gxrnm
WjOyAyPCiLmd6tN6q9f5aK6BSBnJVghK+d8MbO7BCAq6Qb+kqqYhwQwTbMeRXqEtEVH+L+CzV+UG
5HW8hS1Bcc2TsYtYKcSUYx08lSHRer637qY753+LxllzsSMgfjOrsMKgaxuUm3a9ZrfyO0eTIPev
xi5pXbvCaVLS0NvsyFpkYKahHia+oksX9MjWBhLG4ofWSG+qMUzWYDZhX5gTcEJQ9c2xAD5NeGqe
hww3cQsO/9b7AMLyc/x9w0a2Ox7HyDeqqrrZS+xxavfpzcGiO07bc0BphrQ5KSHU0qsQuLV/PdXC
oXd0f4rr6kqfq8M9hRBlrwk4nLHuvkbekXJzqK9zrHO9b0glLh01J2YQH4NzAWPmRWTiON0qztnO
SpXnMzV24ILHpZFwl34Y6CtPGZsF9xhomk4Ao+6wDENWeFA47IS6mtppn+kj4b8lwj0d0tE4uuI5
/J1+P8wIDfJFh2GYciIYPPJLbnt6tO8hNPaSi1wuKT8+bVvdTkeYU1yV1F4IQXuZ+vts6ZsQnWo1
VHTQpHy7m/nTVHEyMxeXQggDpkarSksSIxWw2KuEptXAt58U9SW60g5cSMtprHotkvImfsqtIfqd
a16iIYp7AAioKv3bhd0Zn2SMq5tMwCIrleDE6CzYeoolI+r1EZZcqbD9QZW0fL1pJYwKxP+Rzo9T
nGToykm/y+xEmFz7JXlFxWAuV6Ku8FBK0lnXl3UkIJOf1JzMpKnkhivT84FbFLaj63/8rMTujfTl
6WseLx5bd6rpSivCXMH3N+ISq0V13OR6bRA8H14uw/mhbVtH+oAEsnNWJlF83+TGokOMO8Yl6pxg
lKAHJDlD22QhAAl5SSgZS4m+B3mlKVNQoCXFVO49SZJmw20Ctl8K7kH76f6Vi+Jsypx4AL7dVBgw
wkj2ywbsameHvCeBr1bgdVLNQhQkDbctxPAkyf26dH4NZGJhEbDoXVW8+2Uw65pSo5MtK862/yDT
KsBUb9hbvu+epAiyUycqSvY4w55ixpvhfZDr9tOsJkn8bhpo9lBsXyw0oU3nlQ57uZZ4L5jSsynl
Wf8hL5/bFdauXuMAiR+Io/mhEUtCDB8l8xDbdyNvtI/s6Ri64uxXcXUKlmpHWLczj0k8ei32/kV9
A6rzOLCE1RW7qfjF0tkFWQC3/LBXVHm6qOwsazHAChjqU2LVlxQnSvLWfSg6d0XUk/+DT4MCNbt0
T+zQ4ggreDaTyBkqt2zeOFONgRM2OaW4AH7SOdw2yuyNAeNNZQ2m6p213AhcwOyYV/YU1amMw+fX
5utqftAWlu7Xs90LFNwh66EHCjHQorpFwkDNWPBXcfxlDPcVaxer+0yyk9RiWt5pTly83hF3BsVT
weRM3rP1bUACYUdyhOKnNvtQk0L2PPPIi83z0l5/Hx+nmL4YtgmqUtcKdqCk+1NqmGlpLada/Uy0
v4gmohlRsE/g2ZanG7tlhYzBagSURv7kuiQsciLTwona8mWTUYlOBzcrMoqbmjfBDcmUWJIgMIqN
xUru8frfW5EHig3YqXHpzqof5KKREO0OLRSaGh4p7+xTKZrJNaFuRs14HNgTMgQ2DeLF33fixxmX
sFBg3mDc29jXA3+fRUIVvwen9ztk5qV9Gcdq2oIK91jljarLVjY4ARXX4Y4PzZ38CeGkyHVc3yIl
0kQypZVDbnXksdHjHV8ouDBKN+UPEDrAKlXsOpByt2edTL2V1IoUpmZBNDtlWIR5srvhN5nZ31xW
LJlsCdk2WjY/EsNbi7oQUz2HhAqLDnIEBTOV+qw1QyfLaGhtvIZKogqJkeQ3aotVah0klsx6YiY6
gCdG0+fbmsSMKb4DgTFxdLgb7nXzUmSpzQ7BhfKvZG9aLMWNBMrF37/Rk5nVoMwWYUlQhnBWQaeo
oRIFZ2T0bshSbOPnrvCbZO2Rvtd7ZDjNsVQBbolSqlMeeI/SUF3zZw696w8K71IoK410oOgRY+Yw
vg/80K1vy7Q3DgUQ7hyh/WdfZfR2fEX2RkV3hTTMxf3ermbKf4xr+yuemy8uZlDpy3/1aRBUpSUA
kL/oY95yv5cU41BYiD6K2OranzJa0PY7syHAPpSEcaQmdBDzbPFk9zt33UQ2FA5SqWLjOlIIBrJz
ipEyCoCXVtDXYR0gygk7dFLddet0n7Np1HE6SFL1w9J/oVLzCG58C9f6VaK4bFixYYo0j1pmUqTK
+EluTkU2YeurHBndt8QqGL7oR4A8D9AEm4BBve7J1RR1Bz6OVwmC7IJPnB8Y0ScoZjS2F5375/0W
OrgZJjPc/E3vsHzD9+n35w/y4Tx/1JuaHlIRHSLJiTifdl3URgdOpBwCmnb/zR7TTOds1OjWleDh
ihOGNwosutfsHpra628WPJSsNgs1ivxLc1k5bEyvUysaSOa60YZZ3MeZMAzEycBsi90uDK8UjQtb
iih/W2z4Gl4AVM+oUCTxOSj+GHeff54en14Os8hdg3xWPFR1MHYdNUTRvwDnH+LPc9EtpTWBjsFF
ndlBtqFbD9SXKeeufBguoxgcHQuETrqTCAGjmAw54Yr9KYePdtu0+Lke+S/BLA0Wynj9EgUgLr+f
7NJEiIqTYtrYuZ4ZNoywNKATf+xZt2LN/O7XrrZLGZxw0wGr6lrNcNVNbcIEd7CR81ZJYGqMzFB7
KL0bb+c04s/+TQzX6G1K2dmdhUnfeLyafOFgUSkDp1HhMVrCTILaIVAn6bJuBCtbducZ2yCd9zXZ
u9ozIx3l4U5OvchZRLw/dxXIX5m0EXX3ViVvtA3/fNPRxozwuvEZ/BQ72jGjSm846qWzsCK9rbC6
uRMJUs+oGWto3zoSutx7AnXPg0iNduXfKLsG+AJsorDP0bd6ZKIR+p5Zi8gX/Fs6mV/Rwe58WOIq
5J51WD+tSZFEVyqruy19I4Q2StE+3eEd3K35VYnRTL/dXPh2qalO9ZKsDbMnqjaN26O9J2rOUzPr
psYJgvRzmkDmWQmhh2B1U7ULzyQ5uC0fO4Gk4/S5Ukk62+CbwSTfEjWtBFDYfbTW3TLSnEKh2Hhl
T+Bwrzkd5ixsLHE9kXkYhPiadmqGQkGs8c30x77jsk8/jPllbuyNS0nVo55RRFmpGKa5ZumLKaiF
8pWEJOgglOMg1S92JBSAcr05aaempcgLVGK8ZZct7GeheFjHCHRCR/UyChJGMyxcl86+wAsyzfkX
GrWlVH723YtkfHesv9P0WacPpUCBQXUBPemMc/fTpqzQr9MKkWHpjc0+DXOQ3fs+ClT94uH0cqJF
hUeGp5w3yjVmpCKl6gE/gcwZLyUm+903Fche7ka11CsZljgdTmnVShO5mQmDiLL2DT1rh9vPdz8o
aftuVHpX+9eFc9UTRfVQGiN+jUtrn/VYbVE4ZWbfSt2KvVEnakzYK4P8YPQ29gpPfTOj7TvsmXUe
Dej+DXHh33KWDMBljcGoZYWWbKYo8yTnnqu68QRcCcDJzbY2lxDXHmWOgoQsniAdCnXV+fZYQLsU
mfyFcr+iv4d/qp0Z1Mu+LtAKd2BtIsLQ7TexsTwPGf9c3fiTB1cR2OeuuZZn3cr7T/na1Yw0CmEd
WCn526k38paAs7YgSUHAesuIeR6ZUXhoKTn40/YIXvQG68HpF9ZZE354e/zHEyURTF5vuoUObtIP
nGXF0E38HBK5/jkXCZwvy1Ym43tzEizhNyR8w7g9XKWW5i8bq6+YhmY3VT9f+/rosa/uNYQsGH3a
gpZQaB2OenR7s0EgaHkDxojW4cFfWOmiA0EzGZI3rutcIoNhhFKH5LzWfE+e3rnk2cwbjVu6W9wE
h5NizI8i6rdEbeOAvr3YUW/MxBZBvMpNS6RA1+1I8d5MgmxrHnEs+cW0CLjPYm20QzSuPZOMPYhX
6/nc3ZhrGBo1oESTFTlOMucowX0j0PRB4/+fzbKmmkdFBKZZjPiI911szyUuyFmbt5HjXWfZdUXy
J/Gtqx0IMWpRvibwS4Bsy5nhYh23IbE5mgLni8F9zxtfGMlaplV1mQsMFdYuOdBqk3xliggdDY4J
9PcINE+xFTo6kx5l9he9yq2LhtrItDvJFW7dDLB3shwo9piNL22PahUPG1evSqJ+l+wCU8eoIJw6
tVLY9BVz6EwimgwFmr6PaRXti4zQNGXiS8W7WnViufUtay5r0s+umkqSIo+Kddcm7nrqNYWGF4vR
d6ZUb9HznAgSNoc6UeQlNJMZKrglcb/Z02NOnMMhZYf5nHIRCsa31CHvKZcrU02gBzB7wHwuMFph
lsD7lSsUa9o4gjRX0AzjSSQmj3/qspDzyNf3BhGN4J+Ypku76D/1u5Oe69DPoMRZh0aLn39rZSqz
vftlUlgFf34FEIp7f6p2d4GJH9j94K5UtiTdnIgY+BV8+P6/zGIknCfFrKOVb489zqXy1ztpmrGb
Lv6f5tnWVHSEg7ROKrcNjLAb2ur6mlAkRUG9J5YHNOn/f7FwfMGbICeVK15MfSmqoHfxHRf78FP5
bhB3BshNWmV+2LdGpSpBMuUmaXDamg4etzipAWIkprgKfKMkrXXxkscl5XZRtU4VqFoCE7UbgfDE
Sgl/JHLW82Wxb6OoEVecAZD+aZJOnGgR1aUeCIFR0gbv1KzcOdb+fywHuwZzzmxjVv1mBJ7MVwIe
09Awx6XkRhVfANaFURo3I5jleK+vUAQqOVhB3H1XhlWh/miD3glL4PlevdfEwRD1k8MIImFzyIFI
vsSH3SM5f9o9rZtp1f6FiBiTote47J1ai12Q7Tssdd99fD8ndwQ1Y+Ymjtu/+Ru65rwqO+CxydV5
TbT6msP4vn65l/i5vX61BAjgi47LMTTbOi4u6BxqNPcgbCvy+jNqyCAaKCXRcH4gZ/SPCnPJhKT5
4/ccJI7wPxk/jXxFdDu+ZdhS4Sex9MTnF05S+eWu9yx4Zc19fbFgR3L1f4E5QJSwYxLLBsYGJJu5
R+TvnLCsndeM4FFt5xxzgD9yBrJ00Q4EPPotuWYR0ziuqJLF9+hvxdahqEhirijx3WFLiRuINQL/
J2mg9bSWZhujg5MwzA/jS5Ip69Fz00yX37/25/FHCuIxK/JrnBYYkIhuymk2hH4UFC68EooyVRp5
oE7atkrgb8ElzJaPKzfQh+G46AH31ict2hfvdHLKvV1lgyKmNhQNA1VE47cR8AewhMYE3JudEC5v
5V2SVb2taytQKmsQ9T3eKkrpsQu49uJOsGGDsd4YD/y1safu7/xzZfq1r7GQgLDAGr+Geu0VwNzx
mKlhY970GwmUM8LSK47OAfc2qMrLgLti/VPQXpiLSizNxFlg1YCbECxoV6eg1qcBJSM0Vvwx2OWL
umdat9c4lLbeQkoo/KnOcqC1zA25EsgWYF5KASzdCfVU5jV8TsOvqmRgJdmxQnEcjoT2fn22XuGC
Cvshzp94inS99tLf925NcQKtJkITJTqyBUoWVZsY9bWGQ3j9IhwQ41xav2EG8QA/idTBda8SxQbe
SlB28dgtVaKQ/TSNVbHnmPqW4tsNOofHtbios8RphHWuDhp5IJYGtK6CHXGmPQZchxy/MiaNiY/J
T0x10+3kVcfQbzD5ZrX0dPMQ2KHpQ9ovK5t3GArNWV3cjT8x80H3WoKZR8zXrQ8AGBk+VBbymlZV
0dI5y+V6YTUWD8DcqMMgo8nXd5zJheVLI0yDwl6cQ5PrMT1qkpCUaxui0DUm/JXalgkihBMVa/Vj
hMs0B+KR7lcrTyh5D3kW6TyMWOR6Z/V4Wn0T3uVEJ1wNgbRnGKzJ16qUwzvRtFPpPajLeKXYLj2R
lVYDKQAUCTL/WX9Gl5rrzBT1Hw8NqYsegpcc+oqI7sDXo5xjiWwUP4eZ4K8kU6fsf2liTNoRidY9
2bG7CVcoUhyMjoDJkFhzfEyXtsvyuxbabpqX+M8MIKQC49JGdSJ01UBH0k/mFkLJfAFzFnskTNJD
ZbLP15JQ0nvkuq5KcMuyjfjH++F20Ov6u2oQuAGwoTtv4fKErcHd7hDKIlLQcMtAZIb62vy5qPRK
15UsGpj99m059KM8aycrNw2nMshfPmMmXtsY/VGsKzuJ3+6ZDGVEPKeKscFo4EpAZoHUrMC7JqnI
yvLvCp7hEErO4NEEPitKnTiYqMaIgn0TwwthFzl8OOnlqLHc+K6h37fh/pkyoGSQteH6oL+oQCFt
ON1QX/RVqrfGGD8eGwfJ+uYDtmiA3Eu8zw/a/GRoxw6JGoBQ14HdYW5FtJFfgMSi05EYVMevR1tC
lAAH8sUME1EgHj+uq0sdYQxxgdahKpzWltHq12V3tOcZhNenWvKkzN/0AVx7Mk8rCwudYmgEJs0Z
5K8hkA5hbYlITyokgCMshoXsbqmShjwoYPRoyK2ILe75M16EB07RsRco6nqHu2Q7Bvqsbsa5+Mxo
QsO4Cu1CRnlh9NNFWIfnc7Dni8rkDzPTJcgmgCVEGPxH4XtiZsTbDagdZRhMOkYCpleIRiKPzArX
TgQgn4yFzW4kadneqErtka77gwSG5KBz4MvVlkc0keGjVkGDvuEoGR5pUp7h5IG4S80TOPsEk2gk
KTego2vDHopb9I0A8o4Bdwg58eNdbm08bk9dj/kP6XeLE3ZOk0WFIWimc6fynixbd//IpR/gBy1m
1GT/80NFoVnukfiCIsOotgNRTTCHpMXSfYTtlp7K/Y2mtotVchJurUJdQdF6wg97ygYr40mIsXya
4adH+NUvaONN9LgXJlBsJGrbHpVajiXgUsLZMF0umPzSiwZCqWe9vUThUQEGcsUGN3e9GW9Kqyaf
cppClBYQExlW5isZkQJCoQ7UB144UrN6G5Zoyo8UdVb5cLaMAdSoCAyI6z3SJg3jiMZpT/TRphY/
Ga76ywzUIstwQQnUpub/Q6na5hAk05vOTYaGC2KjyQrODxzcpB3Wnp4LsKLo1OQ/7EjbaR6z8RXT
0v4zabPn6NWlfNz0YZNUfkG4NDOma4E+TdEks8dqvKqyui/UFD0qBr0XFHlBcJ6E5anVTMyJMhVg
n62Ofet3il9Z6CqRSQ+WEuc9OxrgeiAITfWi4r/hW3ueRXQP7nbDZwml29pPPpZshbZcnWc1dWIv
LO5t/IDLiGqZfdOcj42BEXbdmzqm3K7zDXv8FeubuwAuQ3IzlXM6z8sKyegRDczEGmixLCsOHngw
3zl+RDirEn9ho3u/XjX922XAaVpC9RVB0NMC6YTSL4s2dmMuGDNCJeYZ+LqxcBpwT9uubZKSuaKc
3/ejye8bgDiay+ccyLRrPjfHSZgL/hOwY1rIj2Ht1BRrBGy8OXIz773XKXvpmgdd1yNp5tdI2MC3
cgj09j78lSWfy6hREMI/omgd2s7ENjuHw6RDx68Tlro3v6mKEvVCAC0J5h+Oa0duO+7a7V4yRD42
8VmVtO+BKbirz4FwB6NqZeffN8ds+i/2scUoTKNtWlwfDym+23J0WtjXSfsTFZaZUrQUWDjc8Gv5
ttd432QTjpYdmx/ZUJAkL3ivjL9OhyRs+dWaszJ9yHPxltTafbgndVkqzVydwxpv/fSz9k6rBzED
kJI+blaHra4p7dtzOXhP0l6+IDnrO8SYA42REJz0dMtUh1fYDAAZ1UPU6XJzHQU3sHZo75yyTpqD
VljduNwQ+RTacuFe4pS5O6p73EbhqUIAZzaFC2ffQx29BvKvY5wBkNAZxkNZ/sr8K+j8SaYjKifA
nlzxAXwR4/3euw5j0xVWFFNffGZjTINjOhoEwiOt3yNQLICDIDDziVkye4l2ga4zTRi+PJxZhUPg
h9Ky21vkCvTxikhEy/QkYVbTu2TC/AaO7m0NH/yyJEz9opppFPD17z3eZAQKaX5hLXaWwDidfNXC
d/IMquOF/xu7NenVlI50BSSQUuDG6MdbqVR/z6cznLq+58ljszAnK8pQ3V1NCBrDSVrDOzTSEduQ
W+vjkU4u9hwx0VETVWP37do6TUSiCcdygesNRZRgAG6mw4VEedqPAH22qA+OPZzR3FR4i3Vs5yt7
WUZ6vNFyLt6H8+qJ5xEhTlQRCJrAjEcY3n05oN3Hd76WKLFqgMeGoSTZY682OG5j865yygYK7P8L
jBtqogMtVTTKzbV7IINRVPf8CuRD99SzpiEWfJl5sQl71VfjGynEu6BZkrmHhwArQ+ibqWYJcznE
sJGdm1mRuR8TywFtJ5dBX4vVAS6/XY9BLgE6EM+tPQTmK18b/8vcF2S7t49Ere03s5rWl/bmqQ5M
WamsjghraG5QTkFUxWgE52gdgr01uR1gSsFYqNTqrn7ALOsxHyhRdRpWCymxODvtQ4l1L84aLeVB
6/406b59QLkXKFArHGFg2M8k78vjBBeLX1aqQTmx/Gl3jNYTJssGtMdZAuXimnJF3jbfTs1o009x
Q710ywICmNcc2gdnwmIc4ICpeqqYdPHncWVh3sZ4LAchmBFSoQzn1W3OXvWGsJnmiobLCOGv/QKb
LyzHcbmcEbDmBSnKspzsFw7mPhvISKfwJDbzQxt8VnRRfegZ2ctdsHDekAX7j83gRfnWOKiuWZKP
cRaIUv4qWZSRQqNGN7qhd1czvV8i9zBkmue7hImxS+OP3Ew12zt2t3U5F9ztQ15W85GSbxBdz/KE
cd3Ww0y+mwBgiRsyGVF5n1tJFUg12o3ITmCfxV51L8LFTFlCrmmDS8LwxIpkaAjNA6Sws7RYhyTb
goRrNZ0fmhRIBZ+LZPZ2Kdci3tUFj4cjbetz2X1uyVdTGickjYpTyIka9g5DYTM5VlufABSWGuSg
4g+hhB9TXZlVD8WjQBB/cbkw8mh4Qkkuk6nLCIjAG0JrBCwZdcNJx7QByQGHhhDeD/BX3iB6e4rw
i7kBj32uQzuAdfJtCCYNv9z+R/dVa/9fCWDFt0e0/jj6kxxyS3BuUkNrfmBAAfyrllOVfu9GqiH+
Me2qdErEJc9qWzDvBYMSytmSxWgdvj8P1MSqwnxeKKC8tamxP7UaZJaAkYMa6Yg85Uw8D9KzqIIb
vAg0x/AC6iBHw/gUgzJKGVrNL2rpvRE6G1AP2QPV0tl540EIoMlsu9CzasJG20QwyEqqqCvygQ4T
CDe/uiza1KMbE7rRCzhcXbEOm2YuPyZed8cAjhaKm1EsoZs3dGkJofW6ZZStrfpQ+374yJqa5WTs
IlPgKMCg39qtHv1KBPpUqdMDoLVrtQkAHfKlVdhhFE6jSrXcTChQP4XQtq6u8IpCFJ9Ugc5s1uXs
YJ9jW7FcWjZ9LNv4wJ0LgtX+sonwfdF7AtapGrEDkARCpdOdgv5EygDyO4g7Mzny4TMeLQWAeeFk
M4T0p/6bqajAlaYqpHUgGrAcHcU/s25C48hMB9d26XJ1CLvntVwlCvvks/e2r9wFb7snGF93Zxk5
QUWvjnCYCkPYGzbwxygSYzlTFJhM+JakqGQJpEiqXePtwrZZrpKfVTYbwYY4tIiuo3atmM1HJ3eU
NhtlYNf/+VV2Zv5mT/iWPxAQAO+YGgK/rLbaFuucb17QfijmbVNkGpJHwQOF++J9VJ9pggtCH4gB
n9cILAj9oha6QjxzyIWghBT/I/WaYOgqlvga0mfQFyLZZlsZX0GMPmw1Hi8SRuGYASr/ZDaot/K0
ryj/W99TzBVUCnVz2VkXry1/Z7Yvnw2bKCMuyeh+/Vawai5430BxKFyGxse+dEL/7juOwxpxO67O
JQlMaUgwTrdpXcjeHI+7k6k6whyyBzybWQ/+tvj2g+YO/SuuykqikKe3uku8U2gnPY8/hv6uhSBH
ti3NJ9oTdGYy2CW9JlpYUSiCGh20D58esJr8w5r98UnPFBcUd/hdgM+Cl8wJZxNRx1vrXEDbrtkp
ZmOjQo7LRNtN8A19a8ED/jv2UYgNSn/8oRj9+HyYMn2Ld9AZF27wQUDakj8tEDgqi0h4kHvpSkFu
X89wVnW+pA7idvsGS8MGgyfYBbT4VD90VahDvylIiZkK2dsC4qxRPXEqJfdpLdlDn87rSOWn6LRr
tyWEJ/UmUvwDXVNpTxZNyzvyrIRFyH/Onohf6SK4IRndaDCxjrVYkxAqberqBTKbmbR3hv5xSE7G
qGDu8E+vZzu6UAhM6v94HK8/3UJC5luEX8TsC4ZiaEjhYpzCJnxc0KLDNI8tqkUQl/9nuqYcJ0Il
QbF6FtfMeGWAIvVja1HYZDsvi2iypz76ffshpm9HVQKR69HST7By2ATc/DXFp9UeXgFFMgkj5fne
BtgVfDvldFTdIkLViuvr2DsGwD/I2qJMG6cTBgA7ybqg+Oudtww6igndPkPhSBU0Pl8jw6Pyufop
2/FcB0qZu+5h/aaJcgHJC/QXixN0Z5EEIU+LtbLtfghxsZGAZcV5PaAtC55aqkowqP9aoYcbEUKt
XfliKJxDypawDSFV5qBLna/ceLhuiOIdXair+Vz8JsPd67NCJXZJ+yXtD07bDYokhRjymhVc5BM5
g9hbeaYEFwolZ0cZNBOE7uSjyMoceZRHTJkI7GW4kdO+nYdT4wwtSrrA7bgS79RQi/FjO4c+wAUo
eaNuQmysO/jU26fyDhRbIL59hkbTbyd+On3/ZwfINyXCkBtQlMnsquuTnbYFYyvNGofMa1rckFmJ
bSjXaoSU7CTClASxtFgyuu821yk2yx+gkL68E8CArdEILm7BazqXAY8Za3inO4Qgn05uiTd8pTQh
cGIRj1tTsvjeejshK9Hd8ksi4v4SwAM+2Ce/5OURB3dtaQoBKSfSUfl8mJgK+tGOE+ZvBHZSqFZ4
JoHDa2DyNkNY9Ijy/mlgWe7hBpxXCxagffTUs5svKvd+N+gXPywL60Q4ve9g6GKWegwgAQQw2ROB
rIsNjKiH6Dfwr7IZpV2h6VjI4bntL5iGVCcMNBu2F8TMwUHlYJRmLlG+g+Xp1nSTkmzzK2zniQsl
l/i4E7r9XJUPFR/cDs/rUgvBm38eozO7DZYG6frgoUClY9TNgzYUpNxsO+Hy4GjcI7Vn3ibXBg0Q
jx1B3bCGGjS00GSVTqr1F3pGp5FFDhubgPzKyCm9Pffkls3d+3wyOZ8PYFKLa2oTuhEhrFV+OZJc
yei9l/V5hBvfVnCmzHv9oUAzyLPRu8N5ZTe5lBU7c15d/OuFz97BsqxlR3/FIH0cBK/HQh4F7TqL
K5fQaTYp6CqgdLYRwaDn+NRwCjSTx/f7clC+Psdz748+8Evlx0mjAibbidnBuw6MFc52WWHHR4c/
OIbM39WIMxOZjz5TjKzVphRPRapQ8Amdk1veNAX/kZ/iG9LN/J7tw9qA2tL+z87N5OGUBm4A3PZz
5waz0QMp1C17nBVEvd9n0Zk8id+Ke1B/ZGKZVl+qwnLkgm2+QF1rZM21Be2C4/RGwpmSSeVDhVcJ
ndKDlWkrbTeFI2qRj1Q5Qcw0dWnN6yDYydPt8HecZboaP99V9DWr46LNXn8VJR58g5ZUYBxD1199
c/b8C/C4jr8FAMhOkBoGq8pb4vGmaBuD3QiSiGuoF9q5KpTxsutPTz3/FQgesW1ebd0a+cI2pRdd
ARNe71C5i82fP9v4HhLBl067xQDssgNEpTA7xSV/VkYR/xaOjXPdBvOvfn5DX8mnioT/RYKyG+HF
qdwxB/nKfAdiz5lBVZNn7b864ObN8dpXvJeiAGm1qdk6ZNusVK+vvvcFtYiyde9aowjRs59qdVlm
2jdqcZ2GgVB+QmWGDmDa57I3DSrRvQvu08e7034wTFq+9Dtb5qcorTQ2ifIy50tTqR8+pE/u4kaS
CuRIR7svMC8Ol0RV1R6l6p8V9bEvl9Ti7FfT33v3bsQg3zXclOgiDXDC2ZjVQr3lvTPqShDR4HPs
rERcm/UnxVlc2X1+WDCaDIpf88D1MSnPS91J+EW9zp4hCUddn/a5+uPVccWs1LfZq5flCz7nB+hq
ZIDKhBaedCuq0ogt1QuHQCQBftEKf5yOy5hN6aW7o/mhLB5LkEjJ0ypcdac/ns1nSolmunA5ljj4
iQ60ASAE2AmGntLcQqwvFjxOI5vrN5eLREgIUlu0PDiHym2XppLoyZ5u71DZTWsMrbLXne8WL1BB
xznZJvzRG5C0Oyl4S6XsVb9eB5aBZQh9etlDps47OX0UQewBYA+a0thV/9Phc9mANaP3ytSjNE3j
Qx0ksqcaNKubvgeWDFkntaqWyT3SpHCTyhf7OJnt/zhUZXaG1Vl97+WXbuteCZXW4uzXAypPbDP1
87qFE8b8pxRGfIUE+wT3BsbGFx0nv3ycbrzwlNVQS85NTiNVp2KdRIp4p2kfFGHZwnJ6772peEN+
8yOcgCbSdRF2t9GGgHV4b8b7rlOkDAj4u+vBeA6CxRqYbSYzyVH9nm4x+sDlKT6cilRTkatHtDaN
/1cC81k+8+JONZNkTErr6ACYfNVbzj/DXhFCx/gycyAXkOrdE6d9m19tfriwvwhq2W4tKEBQAJ78
6wf3z7rogXZ9BEC5q4OWJFfvjD6vFfFDsn4hB08kit1EXin5G4/W2jQaQp6yjhHfxoTPxaABX2Fq
8zGok7Tuly6jkFe7jYzGlUYsl8pdYOu6W/2qR85EVa6qhxIPdp2QjIWRpHisdvsbDQ3pChVK2Lwr
jvndMmBN0mHWQnmEn/qVCH5Tgz7INThBlliGwPwd0Xp0jbmjfwwCRyQDFZ/ZJZqaTtHK1OXU6rjP
pkz9swRa36QnYPtby2QV5Bbg+roWPwhF2pLlmWKebdfou/dYNWatLN4qJyu44lfO+eJTRdSvzH/k
2HV9f0AllBQtYhghGW4b/0Olm9O0HNbxaO97Jp9vTsCZ7C1CJfLp/vHjWB+S2OIkdpFk+P46bpuI
V7UQi7n7aqAmOtjEjAG5me5ZHSHCSWwj8WlydFvypNO1TpulUa5XgxFbyE5qQvrg7ek07xq9anli
LkD0qOxvoIWjYpqPN8UkUoPTOV75SeIyQduZ2vYAR/YQV2EHff05g/gFijp2gHKZGx8hmULboZou
jk4IRziyg/8t1kiYL+hITh5w0utgAKoWvjPdaUR/9pzq0IiXb5wfIAp/anCnY/rr0/oECEUIQrQt
wqx0QCz+KqnDJsAN8EL82GwUb2mGT/S4Tov5X53Y1dhEe0GgWL6K7zASGdbYQbSQfiRlNqwglLCl
hzD4981x6ypHFOf2OiEjBisRbuagA7C54dftMZv5DGobmqO6m/dOEyfKWXaKuzY4pjt2EYpHQ07m
zhWUKEd41CEMjfUsevvzDTcBdt1PFBxc7Q9/ShnDFgE7eScMjKlu0CF44vuHk/k/eR3rWmGqp5qd
aEEpd46TwJo9nLOUjaIWFDlBk3Xjg791FEkBHGva8QpIY0iT2XU+qcqJsAW/OMP8P7gy1swNcB/C
8BEB2VKcrYBBbInT1fgl/+WMdk6f5hZs4RtIt7fYD8z5973F8if20Tz4Faz9uEP5194GDEQRNiH3
Eply+CuvjLGMDVeiAn4Poac+Yzgo9llJzmP/eZGpesmu0IQd+s5IVM/8E/MgWARUnD85x3fE8caW
tYErjre7+dzSNZJjRQy+6nfELUxnOAfx9mYoXFmZ+p5b6XSqK2yW9YI6D9dCztuVIGhJeNQnjmDb
vmsRWJSNGYMUSgIh0e6UvElFTb15WOVdXuPOaN653L72ym8V8kPsYGnTQQ1LYX0YH9qXORz0osIe
erIVTBo1D4N92sTAUbS5SlmY101c8UEzDLsT1yVDdd/zYg/hgLBCC4RK/+RA/WDvCtCwWkYI2Yj0
rYNnqhbjD2NY85ZTzB1UoaJg/IdFIJGZjbC0753nQiiPC/vQEFn+ZaQ2iuKnq5iKhBvMWBAdBmHN
w8VbHt+I1r1heKzrLDyMPzsV1kRPK+g/Qn3aGZkz5nxJu2X04eP9CChDJ3QBw0yVNgEmomIlKNwO
JReFjxExVZEaGXi9KNVbBPcPojW36jjVO6siYl1ycJ1xQcL6371fTGJVzknWtzlewkmfXo0g5w5d
eILBEfWgWRgO+LhySlR42VAS+t0IqeHoAoXId5ulqWrV53rMFV1XG/IgadTd/ohRM2mOQ4cJJXbb
bgw/GLutDOexYDr+PHPTwGAKuQQoaQVX/2xtmljVHkaKxHKdT7VaHcoB8rRONxFi5OFCSk6zapUV
6xnXSqqVlhUoj02ajgSv/7Ei6yW63T+bbWQgZMxgtoxm7UrHp73nEOG56++mZatavBHz6z1RJ5ZE
0MmZkf4IrL9eoxHnCF7F2JYld95AcBMTUWN1iXNtmRPU2Uo4TrD/lY4Djc7NnvIffg1ixzWo86x6
ZrO0McgJIPt0MOMb+ZVMmzD8Khu33b9OU2rUTBoHJBo4hJaaJWekl9VDssJdFrqGwySmYxHSRUKV
gbZ9VcFn4hCICUpw46rB1daPJ+qDsFK6JOXzgMdlGsvIgq7Q3kgrrZEx/3ryfos575DuXLCfsCT8
1UZFydjeQH2UtBKOXtoZqm6z6Lrdedm3Irg1tqjmuGH36x4FEIcwAosgjZoafqWlXGz639kHkZrg
vf1/wei1GT/i/4ov8AvBVaKhGW1iBskL4e3kRSjmTb2I4uuYFIs2K7K7NoQk79m2XsNCse0RUC5a
Qx+vdZYSXAsKzzB6ISjvoOEUOHPzbh+5RpKiQmosFh0OfQVH+RfDVpqUH9+Seq6/9M6zrvKX9iD3
/vt61jq1HaoJNsr9kh8G1NKSqgblu78Urk5vYdNGVpYbtQn/eue7RZWiIV/+AuV9p1xOGkgz6ogZ
7VoxsKaboz4Z+K3pmFNZndinb3xWzoV8LJD0DV3nQuFwNLhZ4sNOj7E5wG54kslnXIbAhq1NLPUn
x52N3QbK65mWSbhhZuW4IL86jxuq/ET92agGKrDtcFPcn4qhPyGZfKMUc4Mu/8bNfEX/XJvhz4Vm
fpqR7cIMnCzUKTzf4ickuB/PMbtF7KXey6kOyfwmDSigQQhcDRyLFNOxwwzdM1OycXlqAviSwKNX
Ef3DZAWHbZxfyX6xQwP3JwL2M9/D8KuyzGBkcogdUCfm6vA6A0Kuoh/unR+RC2BdyQOVETLF1+C+
dHKL02CTZ/e3nAO6kWKIEsNiVA1rm58YQCGjqFXGwgmaUzBhNsuwQfw8/g38nwM2CgpEN0qHRLoy
fDTOMGsQem50DwqoelaVVed+8a2nDokQyQz1Ksyholks8rIJqcWUfrMRO5QeXtmJRncVUDzKX9LY
CS8TZOEkXfCpJpwpDNZIi6XXDIPyqfy5v06vkfX+h2p+n0b795te5YVq419T8lSV8opevzkh9Ps+
+FkmlaXc7Q6KioEOf8gyFk1tsvYk5i7EQEuSW/hBuVEPBB/+cQ7P9ObfnV+WQzj2gou3T43cxTKM
0OuCgdvivHM35PurK/PZbq6Q3Sf5pMXTYEVDNViNlpyAkM3x2grpdMYnWVxi9mn4m0mBvtxbo6x+
i/qHu8DA1w+pjAjSp3rcNn21o3NE35pwEnuilNw3IqD7f5ErJgotBtePEtqumvNFyi0XpXO17Ylk
/ep5qlU8w/ZiY0Y4vpQfduW5O6nO1dxBPl8UD3uLA6hexDGI3u8Fxhc3cZrIrApes5GFext4ht4R
MD8PJwtrpn8X0C8t+kIXHRRJNn7rJV6zdCN/j0fn2Gq5KXLjeI9nKMnQatXxAKUk+83cVqqY2S26
JV7GmZjD2Q7er9z92lz3aAXQm6uznq4+62++fHaatAn89bVWTpwc32wvPjcGZ3WoZy63stCQ0rpS
bDMLRt/SYBcJkjepFr2icF4jeTeROCZaMFvHaNvr7jv4htOLHv+4zWvk04enkhDcr3oYMaHyngE7
Xi0GFaTNqrrNktswDcfDE6u+OYJJfvuFssaqDbuoRtLmpsLzIp47S8lYt7/9OacjA6WwQAwvhEdk
kuVEWtLa+SnvM1XIrxGnJ30MHbVBxZp/8b/DdhRNHsehzl0tmwdLHBl9uxQ72elVu3jo0uewUmD1
jGM0b35sxbXqby7ynDl0Oy2+ciVu17obqtKafSVimoh7A7ZWHX1STuu8SdJSkRIaJ9ca72HvzWJz
E1mVSRX+iANyb2MG5P3bRHNh2j5Egs0cG0rFGb+uilqeRM8rnMjrsnpdaFgXzrRmP0CUXafXUHKU
sAY5h9P0n0B2/dpOMm57u5ZHRQsNZCyyILWzCziIQcDWmAWlP44i2bSltjdRO5ftxDsK4cWqdXFU
5AAPM0PsoWu1wMG2QDc1kLEvzJm4cGB301EGbcwsSxA5pn05Q9TqWC482i+xQYsLAKTYm2Dhf50e
mhN1fSsZ7UYEL5EJlihSrNge7lSPAhaSIrEKmlk5ssqCGwT1HNkDiUO5rdiRcbvAk6jR8ceDJPBn
sBSohW1EdNXGKUJAH+dgFy/ylu2vmmskYib2UF5kckXZk6k1nCXFhJc65mjXLdww4W2183EdrtpL
SFSd1rmIbfXq3msJvvoU8zGgWux8cX5V2c7z5WOkVVqIRGSVO4ht0qWzPrBppn/KuAQyE8ISxbNn
7iCu683+1sTNXVl64hk+sp7w76mEuLd3OxbO9oeM2lQxv70+gMF2xgRgE6JD+aeymIbUQE4PkVtH
AbeyfUfLVXdbcrW+S5anwQ6DY1MaCbD6V3ijWRRe6G/1vVv3hBM3kV/MJez3JMn5Ubx9dsKa4Ri3
Cs1+kYH1ICR5GrxsIKrkY3SOGpAdV6Ndk5DHvgZVoa/OeWWoFROv2NhFGwxe5+Q5vdi8/5otoIka
n01Szzi6HbsFNotu7kWK0KaWYkPCkMWmaYzvVfE4BXAcOFvEcjrS8WhmCMz9fkYkksH8lYhVfW0J
B9NiFaK72QiwPj5dcdHz7IgojbClOOz+ANUl0OeGahIgE57KNMIVd4JrG/cENLjA5dVcd44temUY
eFxFmd/XhcxnLcLN9vlrfP6DPLe8qOyJw3JNg4LUxkioPuly1r8KyW4J/tMkkWFmDkODL+4n5n04
EWd+D1zbnUi5EUDESjF9s7HXYFi+k9eySvDEHlMGUjjgQlzYiNyUj7l2Sv6pt4iSxgSJgumAi6u4
jQH7kx6wuWaCQLFuYop1PEcxSamrD5zdT4Q6004aBUpsL4l81DaZqpMwTOdMsTL8kqwNKbswm99/
BJflOqJIQ7WgdnptPJG0qCKyV1+juzzW03Rw3x7Ex0hqWHyz/sCEGw2m8k161SNonyIrt3ZOMrxY
OH4i1mLX07As2n6HpLLK6TwBizhS0zL752MrGV40cPNmJHLLM6upzup7nBdUb4iBY+DD3p7DCYps
T61Y8KIfRwZzpySlE/Ok5tRlluEkpjsNvq3PaB8nQmgHNDONM9myB3lJnmRyzy18uLi1BgPjj6Kw
4Svb0Z8SqGc7TR/grwiV0ERST6xMniLpOEqfnbnCG658XbQzapLiWQ+gJInC8HpoxTOVsLzHrfq3
5gXg1qdgM9a7yFoY7+mrsIEFa5gml4j6KvJxIbqCgtQg5isweb831E7MmVf1ff4mtOz1va2czQ3+
2ngH+1N4OXX19LN4THzk08v/zKlDpjHoeJettwMpWu2YEflKR2qNIcqBX4j17Azb4hgwFd/Ov1qs
pOm7mTMpM5OhM2yl5Je//gGlz8SJ/oM9MOepe2W7nDw9qCvXPlo5vgJop8+KXurB/gm9ETgGwDYo
DK1Mjr59JcfF4NSkqmR+fuQz2FZ8GJn1DAZTCM71z/CHEX0J02jeBSmJlhv+o4XcDJP89mnE/Xuj
x+CmHo5D3T1N0g9W9FH7NLsWLiz3MYPxX692EKYWPGxrsg8JsmCYKhdCT1UC9rY/pSGfnfqlCK4B
8NSHXD6tqGJI8OMmmJ9dEu4jWl6GLR+UNci2vj0MiIPRVcnyEHQSO7yIfg3a2PCQOPvxbui1wtrv
6mSc0dYJyAB2UABGbOMhwVqVJ/gvO4vNVg2HAIW0+t2ZMBGRu8kOmYNVtTqWIbIRR5Rf6HklhxdA
9glisom5wJwfHH93Shj3WwWMWBUP6z6VAAZ3LuJWcURoKnN6/F+3Oku+dXA/0fZUi0mL0ZDPv3hu
rTnQqCXc6Pekq+nATX3ZmHm9nDXx/QoFGofXdlNcbK+t5nVApmZMiBug7UtLjcGda5WApf944E1+
jXgJpgXufCIpObglF8iBvdmJYz7Pbg/FSn8o6kjmV/DbeL8vaEmmA9lH6jV8LJY+mLznQjDG9YP3
dQ9KhXMk1Rxe+Zh/Nsg5Tajg0tG+UJ18bJXVYZiiUUvXpNoziFF/DbrUoqV3cue7G7ZrxtwQEano
AecHWHgoGG8S7sCqlvy8krLkgobOZRtLl5Vw72+cAvKDM8TEKtyHbzSIwJcnjioFGgWynR7sS6sG
It+v64hWee4cBCiRyWMeHFryBw7k6DQU8xwhOI3ckwHuf3plUh/30VjN6EMMpt0HMK8guoUyyWK/
ssEvv/3zR2drpiao4LQ1NAPTy9k99up+3C1GgbvB/lZsmc5fV3jyU+IrBvet1ehx6KNkqh7A5C8p
3QRbFFlEdh74vt7Vz4d3xrHvTv9gLCok3u25DpJU5x1ivo3WbPawopMxt3ZgHU1SsD9afZjGUro+
bwg+XiJ2ZqMdZwcw+An6GSeJKNYVhxnE0r4uIALkSpX5bTL9HDGHq9nFOdkLG5lPWI3xnJA/sNM/
sEK+PQvlvToeO7gtSuxkv5RK0KxbqmANHzSwMGzF9cP+S0tWZKZoHZBh2lKP0JYkitlY8U+s42/U
bCr6pjN8XgvwMpotvh+DprIr1Uc2sDT/1DVtaOldoKCyfQwoTCX+li6Bvumn9wGDwHVyf5sUCRVi
wSer5SZqrNtk2kRg9L1W/ZSDqfS82WuGL2lWhiWfPVJTMh2lgFoH4imdWVFkNuL0cBO4YXiQ/HRN
wJ7MUdZfv3x7pzVsCaRnXnsPhxUL3/f2YVOvxc8v4rhwD7BWH9wfBhiYWVZ+saDNDkFg5KVjB3Nr
cZxp9NVlmVETsOKaMo6U/Nrm+vXq7r0wY8lQ1m55breE8hXMujA6b8HR99y34lma8r25AAAiBcfv
vlZGTwj1+vK6LUdHbQCYA0isdy/bqh+A7BR24PT0WQfhBWiyvpy81xRZb/Dr6Vt0aRDvwWsiTxx4
bZcaucWYq6CN5eiUJHgRAs1mDlpJmp03zXJ2cT7XKOSJNMTp/S5b/BsTUMD/o+fmhzjwdAjtq+H8
14CsKNOcUS8Y8kXUOCxOCRzU74dgrJ+DK0OGup6JJrVj/55vza90qTMyVbrDkncHcqpsctZ8NX0w
bZQT1p1BBYItN+63FYdxlPHMvaT28sIjxkuukX4vxo+p4hc/+kYHFH/Umm1z+ysOd3wic7ISTMF3
agNH00W6F1e0hxgDYq9+gI3agHJdIzdw8jbTqirHf/+yCDVvebybewdDII4SWx0e+sm9qDAR5Ong
50A+fNV0t82otUL2gKRxKLl2RfUMRy5+8p5ipGPLsmLweQ9wVelqLQQ3m10Qd1EwhrBIFOQJ0Gnk
Zu4i8d4mFOPkZC7hy1dE3N2Wyadr2QGAdKCS9FYp6OE8L/mCDKorEPgoZLYLeobrPN2qW5GqkGJK
TPXgb2tg+gvHiHV3G3fTNoGfwKMt9JZNyQOnzN/xCpq+K611JTLi0v/TmO82yNlgeRfI0RmhKyxM
73edd0poktblfrlb6vA1cLhBxeViwgBZemLCpN4dM1pCjPPm9H5MCnnmjH/+qdoGV0q5IlJGOmk8
QwEtBWr6ejXBIPBw7vufcrKB+iM9MRYJRORtb2Ejluunuo+9eIkWXyj+eX+uvBwhqluwFhRn9W9e
LkMn1AlkG7MANgwPk4ZwNv7weFEeIIoVQOMWO03IXwjRjFgyPIWWQe8B7jgLo0CZnTYp+YtlKYiv
M0NHNF+VhzRP+8nXvJL3uDIuRZxnMgY9n2mhszI4cehEZSd0/xzLfQrJJy6MjlxrnJ6+vLcu3ThD
jIuA9FBNZEnVM6wgGZ/Hu8qi+FKzwOOfOLHfoYz9Luw4lR6OyGNCRTtcZ7irOOv4Qn4AvhGlZp11
LwYumlMZlN7mWV32V6uvbbiZTbgOwiruolN5ytPAmM/XimXTiocLIFUMkf0KIa8z1FkBrtGYS3u3
l61jzEwnERVh/ehVTNZt1c2WW/NUl4BTBxLLBdWcnYt8b4NNwD8U5WRfo6nJzwzjDHuxLoLJ6sca
n+o7rpsPy8DQbJAoXJihyoJTVVg8ld+NS1T1lhg2R4OzIvcAyKIF29GkjiIy/eKkiyoSRicNEBYk
3VvnR5lpke5VMJobgnekSJR0LsAO1NAckkE3FhaHDA/BT8+gioDQnEjMlahQU9HQP+EOy0F8bJ2k
0IN+pVTFnlKAN7GbB3+Up/dp1QSXCPwo3/nuLych3uTJ56/gMV9K3LNbyrsZeRCFOqNHcQ8sNiGZ
c9Py66NTGkxjX13ZbeGh9KSwy6u9n6UmZamZR5iKwTsyU6jhSgmHYe63ejq4poDqIWslBYHcmzqe
Zju/vQz15tlvdYqvaDPsHQDywYFMIkF/k8qvliuxldpvoFTnVpABrDmmylISrj7cPaitcsJKS5Ru
W6haFdzEKaRItJMVtFUlmOUwqh5Fkbc0rJmHwqN7SNMtvvcScuDshnWBrvR8gh09dFOyvt62xYfx
m61DyHBOkt0KvjAGDxB+z6npkoBqZBXlYmD/eVvHZ07fDqzzurrf7SYl0jUexz+AOUpilyYFo72n
gc4dZ6S63SrOhTtyb9/hKmmkIkmzmoqXNozHDf+QX4MgjATuIne+sfLEU/7HPzIovr+WZZ7PpfOM
MZbxC4cd0bzq6H/I2dEWU4kBFhUeAYDMvfqWtaM/okOKZRHOZC8zp4uRfHSxRo6pOuUX/7IarVEm
sogMmUL5Ouh1oj1GR6C9s5z5DuBxIeY83H2fDGYfYWw6XR/IiNET3dNBmmwNulWJlxTBY0bxXSr2
+a4BuykQNQUgb3od0PxAq+/mBdQsOC4ikpFv1HsNHMR/UjFrL+E+L2e3GfR5CYyweYVKmwP1jH6l
h85r3TazHZ7mVZPTLeicx+KOsMb0TDpYXwuPZwaKFkSV5GULrUMQXBxo4+3Vl1goLMlfkxsJGU5V
K9HTYZAxHQb5VQouiQjgs6UBHaYNXZVMsR9qn2ZMJ6Aozue/kQCHNYxziJJ2RYKux8CtVyf1KCaD
SgsGAQ3U4HH05/BRZLu8/aFV2ljVweVEUZdra954qkin6i5pCECXeqottyw/ZfSqAOLY82t1gv84
GU1EmwUBEkeU58zI1k/hwl9CCnTGUt7xC1hDbUtb4flCK0REjiQRbXif4GiCNUC8sTNrtCCQUkQj
LrxUTeEtfJ7UMjGzoj7QHtFKIwdBx5Kq1mjmdEUqXvYwr25oS8GkFF1/ycYaV1IDTiE9g3WXTgna
+gfX881Ny069uhvCLEyQN/XcYSRg2QCEvUzKNu7mrCCbkrAYQVN83urnZGMQJMDUpwkTxY7DOjet
I74icKi17kTFUKbCYX9Crn8TCfKpTtlfOtsXI0+geOPdpeROUqGlZ/sahsVTIN49RWtryE+xGDjW
1PlVY3TsfGpwLjqy4KdaWNDso+7fFMkMTIxc9Hj/SLZGOR9in99QR3hysE1hpEMbKHkTlpCU1dRX
pDzlT4+oA6Ug1Sh0HT9ne3nYKVqLbO1+zBRO8zSFJ8c3opJR9BH6yxbtbi63rT3uCWkDODfZiM8b
oSTItLjao3DokKCiEgQvqBUctHSuwufjx2bNxlNNx+SgI7BmjqUWMKWpgY+g5olkavSfJfPU/R/g
7GR9p+bWBGOjdq4CIZf+KpN1npC1ZRcRdqMeGCQ9QyprfXVvJCs1gQh9RycLb0tcy90T90SG94l8
abHtCe+Fg5Zr8Uf4Ll5kr4WtDhZKcyBmKf4H+71/I0Qw60eclVSUlxe0Vx/GLYJN7R8QFqsC8LAh
97+w41/XKUpQ3NLXVYuNDU2PdVc+7Oxkac4yHDot7NJLaTicDHxNboulWsGXWUOCDkNhNKHzpF6R
zZxlRAAH+vSwEBVGEAQPWF6iUs/MlEex7m2TWkWtD48dJFq5MuUU4Ni8KQOqmdeSAZcGcs9oEtY5
teCbjcTSw3qtrj0WnJ2E7+9KOPvy5QBob9G0LbN27mwdZODdvzsaBPi4LHzOzv/1HwKcwWN4NjWL
TsYNhroWoy7bov+gIZjBrE+XsHSNi9J+8030akynmoFDifCdY5BaTIyl31s4+JVoeBlr8/HTU/9N
l+f6XXRmsbqU27lbBX5+WVqCJjJHtaG0hwkVLJXtjlVd9Am2WXvMfwCGx4Wv3Z9dewyMGRKG3vEG
zEmHMLrI6aD2AaBFsn6P9oBeGVWGQzqZ/cq4iZlD2zV8IvhDWQkWA98qILmfQIjAOxXXJIE6BAuH
5fPN0X7wmytIwUlYfWY3p++cQbt0Scb1CazoEl1ZKQwXAWuZzvIpnZ4bJdyjbR5YRars/3+X9XyI
4YGlHwWMF3AKiM8rcFLnllf3+jIrzGVNvFE5MImqDi+iSEQAN3DJnJV4wPzGf4KdTiueg6XiTSeA
2qeF6K97T7NqPhGhPvPEwljo84EjHUnrx6mcgmWvhzz0LKSsKHlmOEONYH0nWknQCJVUUBxLZ5iP
YWVA29NuH/lS03FKBgLXdehsMzgB9JHk9WYau+28uq1n+zwoRU8tnMFTlo6L69LSX9Yb50n9zs70
2xCH5xlpI6KScVRm2gFIlmyKbzJnagfg+FDIvk8ZMr26ohAbwJixj5gF+1KzVW0cdfsqpSY2YevG
ehmIFwWT9vRtaFfvVENhvMj/zH7+CGmP8sxUKUiM2w3UMHf4fTJgJWjSwFq9MlfFHNfywxfixBcy
m0GFb8Mqkr5qtW62EZrvy+FSC3LsiR+19E/2XJaALdeTLuVlt7B7JhAlC9RVBwgG6hpDcDUmMt6A
WdqgM1jCJUWyajJ053HClkncxGmaQ9wbPqjYeFoXO7W0exmgI+MuLi5VkMtwgE5LtZKDnYEr9+Lj
sqo3tcqnLsCyOa+G5Hq/C04AcWbYiy9N1cJW7ZBytummS/k5Rld73noxA2U8r9bCZW212MQgzMHl
LTzMqZCJzLhYKuETJg7esyxT/o9QGyIVB+L9YCxZ9KGGdCjBD8doufklPP4iNqB9khzu+ZZSE+vX
QuK0Gx1PtR0+a6o1R6Sk6zh4pDNopmLMemEWUv7tfJTt898mCychv0fRLYtjPyDU86HKqb425qo7
lqe3kVK90eQqIvA2dV24uUftx5I5uqGrKnr/jzwv1+oiIUsNbUyTM+kIeSb0LMKKXVK4ITmklOmI
0ujyawqwFagQ/WMwSlTD4ECOIUXh7v0O8QPbcHyiwW8gUSi28RchzM4/vPy1fYXX96WSEr7CXsHZ
R8qppiEjg6Jm216Db3Y7/8HZNowRArSQT3n81tJeU6K2HblobUHqelAIncqVJFkvCGwlSKNBvRDT
oH8vVBsqaA+H4UTZ0bW4xoGM3VAfsMa4RXCTKus12re/TSK/Xp58ehkdxl5IAiZGv3QV2pBf/3yW
ZaIAnoTPAOHJ8OmaZ35yGqG2PJ7RfhyNdpy4bQ1QD7ztdYrp+eovqtUKUj/rV8CWs9ubUW+Dynzo
VUfzgYY4ab786CXFjoFbbgBIIc1POgKTRBhomQ/2vtcN+ohlTz+/6Z+NptVEiTZYyBCr+m1vVM0r
t8o6SLCFkqtZc+MYjAxdfpwk0e4ylf89702H1uEHTqdOVhtILA8qM8yaAxizgdZ/50StauUcoqfJ
i/Jduj1QQ6r4d9bAb5zaugVfMlB7mFnJ9MckisWz1GLXayGUGOJalX07UaM7I6doOdgBjSNy2/kH
VQ6HACuFvRgOJC86/odsDZkv0JobdLGtZ+Z5CpUgFlBrv3sLuhiQY7W3M67sM0CGtXNEuEkSviTi
xpaMf2rYzATxq5nJTIp6dCLRJcwYB2vW3dm3QmdwQBynEoPLu9jLa21YS40cP624uqLC7ZJonvxK
7xip+qYaReMdjZUw6F8vhVlJfNN49j3oEL7yx78UWoYiExpHN22WK1xStBV6Chus3utTaGrWUdh4
flOHpNUGX7B+ZMNVWFUQycWhnVi2hatqtFgY2V2ZLZvIhkgx6xQfl1VQhgREYVhP6R6JdXASOS5B
NS4rg8EEfR+E0A0G/mkdSFu59ZOzmOArOuVd1xWTdxwoPApsWlUq6h+fVLZtvlEddCHiTJXwBIpR
eUQz46ZqSMm+QnUbZEirvTSk4KQKo1hFSRJDPEmnswhPajF61nDsFGe0LDEsSCJTM2Y7M8OYpXq1
LGF8uQbtNk5pRYR6pNZoW0zjjz7r8zyawa2YiS60KFLrNP752N9H1dm0GhQ2dyv9tPujE/WACu6G
KLw3bbFA+npte+UKWPimirkqlsQLhStfMeICV3ekV/Fidt/fe1Td+JxNCMUSMaGWojnkorCj83UV
afCKP2u7Iw6VEtCPHJviJbK4amze1R5lvE0Th+qQxJ+6WAA2paxsaA6Cm0mJE+3Fs+rRwKmx+DpM
j/FUCrVFnnNhU1YfqXjoiZHedonaZgJR/DzLIUXcwnQcbJLD1DgHoqRUa1DigGIhfTG+xjEYylrz
6jqbuayzCGsYacqpvPAp0qxhPPCaT6NcgpJhiPTZqhPrPjqXpkYXNrCdBbnFJPprRAMHZhpIPvBO
4w4DGvmah1nmvnzt5qkElyFTAQCFnFZOmOw7qokTON5LeGZYTXhXIWTiMSoTKv19qC9jrZOOlcMf
dxpb1No9Zn4yUjI+rUN7MEZZK/7FvmOqhr0fo0+oO3zcRnhinwdsTcUavstfCc4c8SUqHWRVT3Be
3rKCsMl5RMMvN5wGT0O0woHAmdJJsiJ8pqcRYmbjrgoKTzaQReIY2vM305vk0IBMYxXvZRJiufV7
aW9DOcOk8/p+YK0p1h9pu6mpLLfN1ZiZoVmWsBpXT6oNc/pJVs+fE245cSMfnPZ7t9ChYyy4N2A6
9iidC+R/P1/IiM7aT2mXMpCw6fNBzb/zZY4GQyobztDzswaqkVnA61NK/lfQ4VZKPe8p3FsWHs46
UnpLmu2+GA66aJz7v19JiH9ON3D8E8QruWzORxUF8269h142ng4n2UoXNfWnfnSw4y+84P5V2e9N
uwuiHJIFO5lHF2OBXUo4hBhRhf5h2qXkyuNCKHyYfMieA4rGLlXlJdTC450q/SJzkfvItZySm8dV
BYO/hVcX5Gc4K4YQnUuYx3CajvnJ+uA0A8QOLbIudRDyZYMGOw7JwAkx5hjFesxVEPn8rbEuZFyP
D5neUDRmtnYn3EFd+/QtlATPdV0D/j/o6kCMBNRDDF99wgAraoGRu2h4ASdFCGd8f+KbBBuL1IEt
5qmQBdNujaKZAjFtN/+U6kJfozoP6Uh4eRwdcd8oRRGmaZvuqNPLqEcZzlYyc8oBF6Rxs1RgDdpI
emUYDLeJcRyyIGmn0ntOIyvgvJbfDolecR8scefWnNBQMbDR9CuYXFdpJJg2Y7r6DNvcVtu4EybT
iWhlgv454P9BgF1sZ42NeAj4OZfqeDKVqxvLg7+2FmW5civeoNDEHNOT8U8eXqQXvvYN3oNUsOMB
sbUesbNxzpAls2vrX8afTga8UYTK+AGr4mdDOMRPec+3uQwryR+wdGTJdNEeR3vN9ftinJWMKVOn
C49fBqzLpDBff3R1VMZYrWiztmFNHGH348MsnaEQlr7K+yNLrElYeAQs2rpuWWxCSnXjlxF6hhjv
ptlW7bNvTrVfXTogbMPbEkPTytCUIC6cLN67+S6EHoChBoHarHzk0YfE2i8h4TTt+MNXPUDBqSf3
23Rjjnm0LhYVlVDn87pAxwDeZ1IuHgIZ0o43etZHI0CHR5KSXHUQqn7APV7Gt8U53B8ALZZ17tmJ
WXFSXYhfXS2yJzCdablVvH7wjaOHDWBOWCO4Z3EBR1ldkmzddU9kSaT/g6u/KS8ytI3Kq+W6D7tn
LPmRlXaKOs/y99hhHhOUCmiUmseT4b0ecFykq+/g9whNi5Lc+lEto0mRpB0SHA3JNae+x+a229lG
X6awFT0XQJiY99seo8ueZzCJuhNoSM1x5SjkARnMhgmLqVpK/BNzp6dUCzAksfOsD2geC1P2AXFN
AuF92q/Ey6QoKOR/tNYPfBX6t2i7nkj67lPZMdscXQQR0CLOpoO7Lkcbj0fSLR3BoAO/ueb3Q8cB
nJW6GbObRAYWcmjc8wRqx7LoWfZsFSvmmmlh7kZmTJYLny6EbUlr4zv6emuCrCo+RIiAWfHRfe/A
9awi2wjXfU18tw/ZqZ6nVr5PR3DMxVznalObI1UDpTnUG9yMlYnomWl83QGE1M/VMfM9aCrVQ2/y
MQz6Gdiv2dcOhWB8HwuNQA3TPWienq3gASLAN7AZl7eK4bZQSRHYy2Q5s2FCw/1DHIeKOzp1RZ9y
A0SdpaqRnFT/ZkicmdN0AzMANT87SL0BrWPNMWw8T7Z37gJrZ/oUlgH1Ib8EcuPKtwjX5KMJGzTM
pa/phPJmzwSBcfmDRmHFKGCBcwGu/BDclg/HIlGQKkjLOUpG2bktrENpyeRLPGigBGnrWo1nTFjp
Ojeh6kiIwdvRw0BG2UBOzO71q0i/4InvUvaqKNyKmsU4QsTPzNuI68gQATzvUTzmngeswPRDLLWE
phgkeBbb2P0eCVbwO1Ow9YjVGpP6NPEMbHd/X8PluXCMG3ShtISzt7AwjhG4IQqkNFM2k9NLViT9
rSTefDnBnFQV5RIbpzLcCw4Ys7PmoYZ/fRvEhS4aYxgf4k7DfrvGylsa5pEIC1g0NAnMKKPhqtER
ayg50sqEdgWWA3q0LbGOVA2BiHYvfK+iUgX4wDlKpyPnGMWie42c6hIvuQq5JwKX12Fc32s3cTKN
x+yApXNx1Bb3O+lXvhtcjBuB0RGOrUtCxOt2HnVmazLO6EZOI6F7FbRr7YliST0pqNXceTHnbeqb
Aj7ULJMy9W4RqBfrHXuP5ONPl2OEyrqh2VoHFkJBx6YUoa1AB105G810RPSSl7BdUeprDiBWTjYH
0IQqrFYuoDZdxYcSZdzYBF1IfTt9B+74FDC2T9Ige7AOIczI3Ez8OefZbIxd6emzKxNA79gONw9T
Rg0LKmWITSn0cOM0mqJYAhGIaBXqLAo/PYsV2hNDtFIi+oFwY0WU0XEsLyPoUggBIfw1crjLW/4O
J4xM7A9Fo2y/frdLnn3waPsLu7vxXerULGIvdsa9KIv2+jePW+TM7EswtcXZe1ejLHWpYZLBBqnb
wsz/5+kbMK7iWAyP8wPGbrkea3EAvoHD2Jak2Mv1FqTwVpBDbVHpeXGICKMq3I8NDeiKeTJt1NGg
7Q7n/BMJ7Yom7mdC8/Klyk8aMVdbjBMIfLa/R0R4z92qXgTdRNNpLOd0msD4b2PZOU1g9iIeQG6K
08vfdqbjPU5ULQfsT54biHupkYIgTQS8Faldz4++k1QX+NSLxj8fRLqlXWdviA2YuBbLj2aR7vJ0
mv7qgMV881PygDkUCiGaFobWpR4rd+XI9dsbMcBX+OX3+cp4UHLiK+s3kzmywtuebWseetbAODkd
nuOHibrBI+dt7qyVDhOmgsTSOeUaY5Puwo7cUcCxU/eUI6Dd5gEc1eaqYvVAD72uXL6m5mYk6jod
9PLGXKeGBugpf3WxVXjpvmTQ+fmJ7WD2J97LjghWFmQop/hNuu2TMaogu0cY9DaFgMN7NZN/9wdq
suMYn/YMSOa5up/3rtD+mqYer/wprlGOE0JJjbOZX9TrB37CGKeB0uvNnkz1kMx1o4zjpRfSqWgL
AweSvFy/XmU+fbQWTIylzJUZ9iPtdOJfyuKNpTqzchK8Tp3FO3IPZz40tZOLaoy0UN+5nPW8LF9a
KQHIvyNlnrzHUL50O3EZFOMuQPbuTE9irgxSaWqVAI7rOb3/HMvKFP2tqFIUeVXWxs1RM21Ivh16
1ESuRQlNmaOdCpwnF28cX2PxOoXJO+5F1ulRURlTvGmlPbDRdjNTXm74SjYuT5Z4aS85s3XLYZzU
a34RkywxsDGrEPdTGt8VAL0oq8CO8T47Ia2KQoREp8Zn/5CD8CjifPJTYNnURxb4vYgQL33Bq0Rw
zyAPbwbWz1YfaxC4L8VXF8QrBp90Rac7tByBmOFQHcBl81eSSs4vo0NA2CHRwrHx/+9numCB2XC4
pIKF/Rw38kMGMCXrwJQhwf/pp5lyhiOJBfSGEMjS5NRrqkcG0sByF0xlgu9hyPELoElAr+2LJHRR
l5opu++Gj9Sn5ygS3JEJ/SHMWoJWd63Z5bwSi6Hp1EP7dEudevjHCAv89xJBVGv3eu0DRXHAhBIS
S4AeL4wfLi+GON7m+YRqGfNgEyyXrrwPx4k90uPmEs31JJXNKIhUpwl46MNvIjdUh/M9FehPJqiG
8wflCxK1Ex1umcZ41rJGYA097VgSzNY5Ht/RUrFH23zCkgrBQ4BhWjGaSd2S5wrBrCRf+nrcMMN4
asEuwrF0rAyWnhahyJHtDwDUoKcusIxHE+CVLsulTcAGy8qjHVmSF169WPotEy8KxBX7SP/qb6J6
ObL9NxKDMvalHCdMSJScDyayBVTgto2inj/11Wnd4ikx+Pjlv0Sv7R+o3I5PBoht4F/qXUVWzr3l
MWQj3LkANPvTtgslknK6XxLhgW4AIm/rbslJSAzrjGjwqb8fXGNXLxLIWbuXq0jEWoVIEV7U1JRO
dRib6/ShGaj7vIXX3o5TnuQyv1zCaSff/JigkqtM2UOGZCeQjoc1HpENQcP8pvt6GnNh7wi6bcYB
x1scfRuxH7extAB6ODsNk5a+j/B+Cb99j1wg+D3Vwb0nyx9k/7pkrz9gbSVW1yFg33n2z5qReVn/
C3Qf5Lex2OI1hPS75ijhKD8MROBKk3YEjQCiaglhx8eMgcyBW05Rghob+RucKgV630okv2jT89n9
uDqKpKcBhjOp3H31pl9fxwsk3zFJBCobAwE07NNLI+5NVUyroVqFSzACTS7GMYt4rs/vbzwKQ4Ve
qZ0SCyLsmllk8729nsMP0ELMO73tifUx21o2+F1wyHR+zCypin28nx3Qhs+1o15DIsla3ZUmFgA1
PSZOwq7R3t6nb5ripmumf+5sSAl7CirCSseoVAkyX7YPMC62tqmi/36r5TnlqcWE17NvZfaqd2A/
Y3Cq3/y3QOOF4f7Zs5m2kNdnjy4NBur85d1GTlJz8l/ukk9BGBrgYRJh5CNN0NP5LX+A4xp5Dwy/
lunaG/YCPTervv4i95Jx+5O6zpAxvfe+bWoJpHlY6grbokmfO9/5oWhxywX8WPaXJh+5cJWxz0mW
wGk/bS2zC2zPwi+lGaNO19ZXjCoUC47VL6z4fABPdDn8xMg7OlL+xhG3qxdKiDN0LIwLOP2AMIan
Bi2enD2vV4KFhSgyx91tf8xqBrRv+69BPDK+bhIbVG5Toqbq2wFnEeFdvtZXVIzP/vXDMk4A6CY1
eSMcUa3dUlv5y5QMgvsGQ7MTLiz3a1C6itAt+KsGWRiUwhqBDMRCn5vKL+uikMuq0Oh79U8srgf3
CMIX48lUtmpeYhamQGRlXsmSrEztLFeC9EpJhc2oSL8E26pEHxvE9UGCW64W2YV9Ej2ITloMm3d4
RpuIP76zqFeUXS92rAmHu0v3zYBIpBR6eOi23minafbxa1m8vv9j5Z4tKznqTIQXuy7KxnZ6nDsV
j9rtBBzl+vU/ZDCXw3nL1sa1so+hd5eDpNIdjdvpkUTeRuhAkQteT4hVkc6M8ksihPt2bfxS2IBm
F3sIGCWXpIveF8SobT88xvXFzUk4E8xRMzQ9IPkFSf2T+Gd32K+7mS2+aLEWu4AgvX+74hF5HcZ9
b0gydzJGN3zKcZ5UrSLJn2XHZ9ZqVT+qHt8oKUkHp45tCH9nyqN0PLB1tBO6Dz7el8HdtY4wq0PD
hVKhGEw/qp70nuADGagZuBQAlJfbitoHtxIMlDBMwGcEGbjWzWv02npaXxXAum5mAFVBLH5sC9+d
3qoyAeiRWkXHLVNewLttr0rceCoAyO3oE3O3YztwvtVVtdd5oJ7cEHNcWAkhEmCzQy5FxjfE9bkz
3x7rXGso8qLG175GI0KDrNp64eBx4rlWYnPzFp6yD7VTpi70XlowgSDvsZPHlIAoYW3L5Axs1wbI
dNuSiuXHyeX6o3fDtoSr4pEMnCzZabrKaW7tzBt3G4ID2cjMxxYpzs+qTYhQvO2xHOpBXki7VBZi
YfHPvDq888b3SiJSCIfMSOuFqnMmsPo0zAC3ZgCktNTa3qgFg/m5qkDqFqT8hkKLIYRislJ8uik5
m9E7zjywNxk5Qw8yQV6YNk3mFQkkbh6RtPV3vGscO13sdpd8nuIIhJeny22RDp83FqaoQjo6vGzq
cYCR5AR1KQlS5T6o4ErWXLhUOPSgg24WHPWO2s+mTqPtMuWCXtHnXxgxiLxJ3b4167D6Q53A30Uf
olX5O9tKsq2T1OEHZmyWf+UewQ+/mVFvsHIFv8viwHloxqUSbEMhG8424PKs7wv/+3gALjaTzN7N
7ZsVRtJ9qSgNloGFedRRtbY6Y4yuJwqoLbQj8HfFwGHKjJTdpArYg3xSkQctZ6eBsmr5cdhkdmGx
1j5kTEIZ1ADex66fpAG2qpP7GdpUc5EJZaO/OsJbyEr19VOXyzXavVC74pPRnRHcJLYlFOpjBvqE
WLle0BqjMUhJCxw04bKyKk+ZhONz0TnxtM/6JxZ1IWxozyew5ek+PkekpFE1BIafMdsFxI/qjmh0
5HQThiw3EAFSqioM1mNrZM4OPk46vhNcPh9Hq/r8lkN4AhtWqC/ikZMcYu1Alg7NZyOojf4uBTrf
JmxPtAjcz9NQrjfD3UG4jAHdZzoDU83NCCrY8IfuBg3CNCisHLJc+3Pf9EwhPID7dQlsNbQ1dm0B
gNgEYY3d5f1iOkAUxGsuMbae45wMWoenbSsQ2Vn9gB4BydQBNl3Cy5Rx8aSIxS0E8YUj+azK3Cka
ln+Ae4zEYI5H5gWv9a9rPwsTZSvzGyLI56dgVDBemdZPyOSBlYvwcOrclIfXns0m0PZSKWVT+0i8
ZUmf1feadjF95aftCUwf/Z2B1VsijEK0wrZbVYIGzkV7LenJPIQe19fDUoNavKF3paF8iXFre+h3
4P2id+GnJX1zTX/YuLCTnk9NHAKzmRS+hPZDPV2FvFN653+tYod2dBqCn0CWuaqLud27iWLwdG8J
ve1bif8qplOVynSQVXpvKAGU/fhfCLlYWP1Mc/MnNrM/QALF2q3xPvj9XeKrcAExE1mGIQlpI8PN
1dUM+ZBJy5N/LRM9Q6/idZWd0uBsfCF5PbBxxMkNEpBPosacW3YbYfyzhLxUPHIMsfqbiV/oWXx6
bsAKQosNG9EVyXp4F7RESbziycftbAg/jBm1IHMKpjIIPQjIMuC5Lce6iR3651kZXIx5AncuGBzH
9epTxWoQqDukYcxg/rhvRMlSlI14juNved2Lx3BW5XGs0at+4/zFDcDsSuTPaQNEgBF1frI2iwm0
Tfqz08DzUEVH4oTfD596KW02Zy9ERfXmnugtAYIEp1thNBtpfLxKTpnlrW3Vy/TinkC8K1aQtlBi
Y0YJ/7/BhdHeqGxndeHdFTwE/VNmjwIbCcnz4x1thZiMHxthzRA4jftoTADy82Oa44DHe9GGQXAj
9xrJHNmAZwhdSZKmisw7nnjpbPbgDB7Q0Y6ZQP4yrevcVgxW9WY5brWvj224fKFJipABmpjtRFml
BuQ28wtnzQZt0XL3IFG9E9sUdBt9RE4KPn9fhf36MpsQXfJOrsxIYjjI6mGyIzaFR34Kwt5S6ETx
FCzEsYv17NL/JmJIaou1PSRAYYCwJ4urtBwQkSLM6jZt9cwE99cG3eU53v1GuWyBhiHngL8shL9o
1A6Z3JZkKfvaya7Zkwo1qhRXCTbaSqwPD1yY10txAwuj0XWyvDPCezdB84ZGH/KtFqelwdKeEMv2
kWN6NuVFgmX2JJAHZ4/aq11/rSHr7hpvCY1pA1wkOllfOMdPIZLm8cN+UUbWxZqalyegMx9oRl/+
BNE6k4vIQr60oix2tOPQVkr0KwYuqMWUtc4MSJaIOnW7E7lUYP2F6lQf3jkuj4PcY8f0xzqJMjST
yuSP9mBC76hfo78nU5y/BR73HV75WD5FTYaj66wafd5ck+9aZdGaeEsqLtVDkg1lJ/Bfl0r5V2tp
R9XPWO0tsxggzvH0iHlGhY6x22rrLJ25w9AqljeC0huA2G1qHnF49hkaTnpD8NWFKyDJBTOIkT6c
Li5jQjHd1MOzttjYxkEwT6sKJd8PsPUz2jksXDstwJ62OWCSUTA+eO1QCGVmd7WA25vQYaA/nWHN
X1t7txdUT08rDbS0iRbyVqu75ynaXZKekbR9O9GNywZD01V6sNx1BARn0zHJWhCM7kwTXpOJzUbS
cNikI4Gzn/fGu7tMVo4hG33J5RaE2qN1/37ggtrup0jutq9FQa0T9k/qnZe2D/3PBoQTK5j0nO1j
2GNA0Gj7TKo89SlmBSA1BaAdJnm0QoIsjxl1L+SgsxEX9HyR+BRym6PXD8bsMx8M228ta9uwPnEA
VNt835hsrG6VNYrGq+jYD5U1SrZRgFmW5e1Ge9TPuSsVWhgP63AUholqLlW0SYO2Bcg1RzmTuj5f
YMlYJA/ivfy+JFGVcFqFujHImLw3ja0MIhfKlikuDFa2y9pOVioB0vTy9EdffQqqtY+p238DV6PM
z3/8q6etsLlkP9t66NkY/V7rVQl+jIB+oN8f7vQpmh1VGmQ8D9RpyqT0yGNHMBsrSq/g1UBJo/o1
6lUfzqtx3ed3at9qUxY+U58EuXz2kg9w6dAbrHZjZmO35NRP+bDHY9LJrnHhomtxrsRuaK9qSsig
x7jr8BnnXBbRg2ew2n+VNLrMsEPMcWT9GV9g+1QQwGwiqI5/cPQSPlshIkEplMyxOqYnfyQnzYi8
ef2aUjg6MNHPIUjErlrFGmtRI+ANNg/6PcVV1bt0MOL/8X9miz2RsGLDzLpCgMKgzvQFy9o2d5GS
nf7knoU0ky/tN+bWTc/Nel3LvivDvuJPu4o7u01Y9jjdTbVYJnFkzFWByQS6BmQVp8vcZXfePMju
q+Byzq8WKUC+cAOby+2AKdcBN0cbve6UhgT31WRTClnh9xOk4BTKJ50XvEHsVb1E2izHBpJJQ80f
THtCqmDxgbIfgDdycuh5/xLHrFT43gQSn17X7ecm/pRG38RLPC8/vS1uv+3h1WMjc24X5TrP57uy
CizEJ8ap+eepOwkGYecRVTtrtsZE8+i3K5brzqtwzHRUJNHlNNodRFIi8hdvDN006tmYS3/teFB7
jYME+8YrqST8tHLQfqTpYrIKklIyLkSrnD3XyOt6nlvmCobIqjcqZStrOzXs9Wbf9tTiIKPDNzBI
uzv7UPAmmYFFCqY881k+PqxdJIayZuauv+2cXhrp/0THVP7c5Wa/lSBd3p6T3uVb+iDJL45Sd2oT
anR4LLyhObHPy/D910UcPzsEt+Vvt6TPEs93SDwpqIV9JG3C6WmcVfL3qehe3WllNjzLPFqhT+Jb
BXBOEi7e7uohZzvXRNWunaw6+z593Klp25AGyfboYs97ILt1gW3aiUqlfyPAuwW6j8QxvAtEGjRs
4WYk7MeNSha7riUv39WRe6MI8spRQpVwndArfS0NrmmaLuT7ai1fypNWZ6ejvWezlVPHrnPkvaLV
LtTCQ6lCfYz/NxqoplhBd9mqZ9SLu3aWNPF1BIzWS0ahKxkXOrZ71bH4CwuguHTW8lZzwOLBdFFI
GIWJI6wYKpnL9yx4GtaXsaTsAS/+fVqkZLZ0dc+PQ3h3bhpujvYTs156ARvyftyOgbRJ3l088vTh
IaE8++fe4nBy/16/So2PggzEz2CEGzMH3GNLx0sfpc4JD7I0FOQmvjwLKW9lJki+z+FKlLHaJf42
um1ojn23Lwaj9Hh38x1QZvYE5/PAn5w/JuaKJKdIBQtYy3gcY02VOT34p8Of2iNOa2VDna4rgjkD
IqoXByI2DGLuuHXRHct6AOEFpV5THNSLpg0J8vLz5EvUHagYfYFQ3QscIDwLh2Z8iZlndDXSrjXa
fHnhVzWOVF/CpJzTj9hC9I9h+hELAtcJxymLH4tstWJqJ7azkTmrUjrO3WSBdHk78/2wT/Q8mSGX
Bc0bGeaNEA+lThuGlMJtpH2AN1q1gFM48fQilo60HfCYhSAIhmJRKI15Xpxktbo7p0IboO5embVe
edYJZD4rPqkEkmsaj9qM3VqAeyDI8TFl7RvpgxgduB//Bnt0/hYNlSfRZBq17NmDbq5LWXnyU9nz
WKDsvzxm9R3K2WByfLTCbkMtuBn7TALVDe40UVHdfuTNS7r73bIReFTS+hTCV/d1nE4s1TrB2FKC
ffpsYOa8ZfO9m3TRCaON36CWtRfY8vvrkyGuaLrZrxbJ3PCAkDPbOnobUdr/pbxy0to7cPJyXRjH
q/T8Jkvr9SAyzwOM5skBGI4k0VrVGYN5ynyxuV6gAB3Beuli5Iz0XBFlkpNmQm/h9dm/QecOuGXv
QIzKH2ttjl/cLkNFQ8Si9VO3JAlXVj5icvgx07aRPB3X4undierinHbRQIyaIQaDd5HyMbj15wYW
GS+vaqgeKCanBmiRbp9Ifix7E6wYm8QaDvHT4JknczPvG2am5TMFcZ2lK7taLDtDfFlzmUcxe/CM
2QO3DGNBj+3r1Cv7fFwERRt+R8tql16CxtDhWxlLzCrmpDU63XbMdA7lal+vF6wiTamNUdNTSUnu
J8OM81UzgipXxMfK378fC0uF6DCG7zdghtT8YDxPadUPU/05fgLsj95S4cVCW6Jqajmmd17Gt7S0
T47To0c0azIxF1FTL3cklZjMNXXbri4Wj4sYfQcf0m1DjAqCWJ3wGnsCmg6v4m6z805FXB1uTciF
aHz+89OR3wQ0ygyngpvvR66UpM/0l6wTxJVk1n2VpKXIjvZ5hVZfs539bKRfi0sFlLgwBa/tK8UC
3CoPSr8ISZVPAsWY+t35KvDQnx4CSpmPdh8b1q8qXKWB44z+6bfkehlSbcfhcit0LZU2EVyJFQ3m
GGI5lTffJ4QrgMRqAmJpd9UdwGvs5DtWn3Px2N6mSE2sgluwsgCWtKhFJnUrmes2g/7vtz9m9bpd
rAJDCMr+cTzr/k6nP9JOYHQwhNZ4hFYFoxyHaFS/d9xk1b4WNjq9gw2XrpARc9n4CgujQ4H+K6WG
8ZIcxWud/iovC508v//Q9pvE515GTK3XfCYkbuZxMGH/lOYQTwxjvoDg3p8B71ibvOmEqpRd02Hh
iplHuWQEckhxdEsdK9K1+B+7VQMAvOJ9NsemjZMjHC4bpCeuvENxquVRNTsMSPutX+4qFjYb38B+
6wA/thIYkXugOAmX226aELtOH8nylgeYBfscqF9nma3m8oH4RZZpzdRUXjgo+Y+tspv165F42F+t
9NL846vVyNmWfCN2V+7ADRtXTSIbhCewLhantYnnSFQOp1P9gQ4i/hwzkfxK8fzbhYpQHoRUhQgy
MYMGHJxILzPIsUc0Pqfo+eWDyksFElVBIQX4pHdU0G7NuC6z4WtHnDN8rMMcBJyG73hgbFeZQ1VO
T9Im3qSf0T8ws9oikcaZ7hWklIgJ5Qapsp+ImgCjFz5LS6HLU9BhtddlCyXTDI6nSxEFuxH5LFE6
AyGo22Z9m7El06vs3x1hmDTvS302i18X7DDIucHPGwKBsIZGe1jJkFS9YYk0VKpr8MGFnJ2rOUlt
Ui5jOVBFmbUDpEfYY9ZQZeBRVIR0r5tba6FcvgDyLTLrSov/z5QCrxC2GNzo21LeNp/yGSFuzldR
tEoW5rBBgm7tnkIBrx69RDNJzZC4N6DNdCk/MXLDMXH7nzxlflXEaV1N1epYvg5/6ndLN/g3FkVk
VDsMlUt6lKofgfi3k6WDFVNMJe7lLbtFyliww4LTlv/MWUkqpOaLyh+mAl/wbPOnYPQ+b2VkrPSb
/ew37RrBzh4qTUc44/JWfzXkJveHztwidusLFCJjVLqZ1OlKXFbrDO8ld+cCh1P4GK/mq4xgcBCi
ezPlmQtQ3xJYcqIsb0urDT2x9VACgAh7q7e6RFu4A7ByOpBpQRueBScxb+zpoVITMwVXBNwhgM4S
7/jw6XE8BfqeEnQJyNmFxTrBAsrxRcHeyRxUg6rdOpQvF+4y4mlKJYaYYs9UXFJ8mN3/x9xhFyXX
SvrvCoQ2gxx6AdZEulx9lBWG4ErAzPsK7tXCvLfdXwE7yqY2d7ik9yj9lKUSNpN9/iQItA0YR0Cq
4byTTIgmsZK8+CbPH6ZEg2+X/7xfr0uurTNXjRa9eiw6pCz3KczkwIj6XEJdezkQmEMkweS2WfoL
FDoKDLImiuJmJ6b13/9d71T+6nthidNbaAGWiR7AOnkTS/pcmSVU4rJUS2V82AP80L2WyGiKbpKt
WFVDLT/jk15YkWnDH1aG6N+x46W6djoFxXIsUXvcGe1maD5QuSzdAqrWHaed1WlSWBXoj7l3Szn6
hSn3iM3SLRuMv1d2uSmKkqKVraX0EsT8MX7yGwFs7OQA1C4iSQO5NguuPMjknD9oKPF8tdF6H2Sh
wgN8mvnypYf0sQ6cLjxnB0bZAe0DziJfkjNC1ujzOkw5KJUGNQGtcRd+t+qwKAEMbLTjJJ2XrmWA
amA7BHglIzZ+pk2BrmF8nltNViHnuTEPOrNQ754/mpoyvT8NVlaMc6fRmgylp5krHO/MPARZd7yq
BmX2cnG9qrneYkwXZS+ryVDXQqdS8ODokIzqmoiIZb0+Kkkf7ojcAafMtyIHhRCkfxnOZ/Zb6OsU
zq/7ubU1uxlrFj6cXhtAhPpgz5Bdq/ZErq8JQyJYb/CdaMwsvY0qhH/n1N3zB2PDCj6YSj4NBqgr
3f6jBRa7SOr2qZvjbfsWi9YLkuZbM66iGcZQmdRkUYoNWjkKIQcaDcBgRGKY2s59SDQuQN/NeT53
UnWDGflbSJTg5OG/WHVWcq0nZmhb1uq7q4ThqfM8RnU0Addt8idc8uFB4/o1ez4LjJba+EX4PziN
FepulbJnOBSJ4QP53O4DZ81T1LY4UWNveL7kExF8bXVG0On1QcNdiYzUivlfgAxK8q0+fpSTg1XW
4XNYqHHx0wrMMWKndK4fEbuiYrBGgE5aPsBNYG2h9I7E2dfof/1z0PynfifeS3TyO+6Dy5NidR2A
asqR5JUm9VhnjCAi3xWsOQfisArSW/1OJLPJuZkhrMHdvgRBXk7/suNhzY2hnZQk68hKrf/L2uZI
XHv9q2Vapl3SECW7F4jMqN95FHM0DUVAnLlFZ74RBNOdEP2l3ueGu7U20+s+nDiO6bLhILjcs4c3
imqPeEV+YDoTM+LQVvoGOQ2CdLyt6ROY67Jm3YmrNoVqb0+9P+MyEKTkaiQ+QR2lFkwXlOU+1ytl
fZ8QNjhIyw6ys5Pge01tHuv/fbftcRxLU4WrxU823YcSZGMno1hYoFEi3JcyOy2PP4Q8J9IOAjOV
Jcf+ein34qpXxT1Gvfokz3efFxFi3YvqjLf/huAJuR58rWRifB0XXWqt9SI9JcrEfYwcJoDAQ22s
LY+8tJLQqlk8aLYSQT7/hzs08o9cTXo74zRioDueNb/qtc/zIL4y4q3jG/Mxe7c8/dMLwLqqIQQa
0Zr6VrtFeM57WBhHPBeI/kN7sMseGGVS16BZwmlb1vkKqw21xIXq8cxSHiBLodcfMrnIErwR/l/K
co//4yERmwBNbYfrAYz6zWGvqcnAUDmTgGhxTqoSLiGJMeWgh3l5GVmnZo4cacPr2vjfmYE37Qls
/qIYjoWly8jbw7HASD53HHzd+HISXol39vGoN5ucGwQUxAYE+fetDhZZIqlMgLDXLJ9TQO6/m4pJ
Dxok4c7qvGy0szPG1++K7wL30ZI9kVI2q/nPVq5Ph5LtR2m4/QmmmQfJeHQxtuVf03s+HQAOAfLn
rNEHbB5DfDN5toiWByg147+NejwtN6z0axCDvPH2qQhGUifbxrvwo6DO/p8FbH1ccL3GWVs2WUIe
NtS0wLe2iYDUVvzPYVKvji30jl8ulN3934/dYwhzgpPHDxLPcODY1OhrxGrk29nIBfIrkLNuLwLi
atBnb43zsMuvPMw+6TPCs2V+Ptj4DA5NzBSOqDtNfBYG6569jGsGdUdJx3yQTBuUB12iQw6ipbOy
oEs4aFvxKY4GCqggsg/arOQ1DJUaAEsExHiOOvdYQPOnuqneCnUhLeaAbT32Hqk8ydY78+np+N4G
kYJn5VSnuxg9KCABz+3VQYWzpYd/geagsiaw9r2iJK+7i2vvnaV/Mv2XtCoRy9es8W9oZPgfUfUq
XUtiWS7Hs3QFUIIUeO5YIdrXColOEQfZ7NhnamG8SwKAKxOGmLMxu118sG3Bq2L8SzsSn+LVZLHE
lIwn5t7t1j3LP0Kicb0uZ+KGrcUIrqnKJPuIxp0rVMU3HiKAAXwwqVA1tQBDjluWO//MVO1QIbrw
BZJIG4euEM3ONva2ix9T98nUAlKv7fB+ayxcjrpMbqnc7PziRi2XJpY7xaKznrZeEciOwh4CJ2Oc
+8z+VfWxCb81/7M2PQWrEkTStcMEi929N5RiOMS+k388bmpcVG5eelXwG+8gLno/2T/pqGJdHSRb
a2QKQOCDxKxwh9Oc47RLrsc4sqHbkBvNWJB+x3km7/3Na1WBkN/YCGmpJOEILarz7vH6d/X5GyEz
4lkgEx91WSIfrrYXpsxloylcZQAbIapWdHCMtKdVz0u+XNaOc8JVEuvDA3tSWmQPSB6aBSKmOsSr
7su2rEHAFvToRhVIjmNZly8B2daAr9Js/8SAwakAg0xVNOmH7qaAwlksrzPRwzPRTgHVexv2jF3U
61UAP98t8VRc8C2BaaKsCBh5yh2DRPBFca7Zl93oTmu86RRtv5g0K7iCvu3qvBd+Jhg03EIHfVRb
tWSPIYopgOabVvei0SevRsXw4mg6RjN7AmsChm4D9kbY+IZqDmXu03dMB6yAMeLhRPmp/83SZb+l
TkhRE8auQsxhpyom7edptszBA6O5/Z4il3TyuxQK5biTaUraVHnzjLK5zJOI4jA4TZu6gg6QkIUT
BEv79Qk1bvQVq4VCvQXyo90YEjSXfSEIG8EzryMWsdV5oOfz3d7ei4bSvPDdVMOWKRBaT17S7fgu
e09dw0Djcz4GYl9UcuZfTFfOhTCa9sclX8RQ6ba99lwSgNvSRuMSaQDgP+nSSBWJjl0QqaP/+c0E
wvY1eCQjvptLHUTnoQpz4MvfUzLKu6eT92yEx3huvrDTp1qaklwHEHaLWDoVW8JCS17l4IhSf33+
3vZlKFFXPU6ICWsa/n6G5udG2Bl/OjdHxI2MlW6W+Mu80xUD6t5oaekl/PKX/5OmW0F8Pfn9nDaP
sOVz3LZYS3WZ54ACFMrc7csEvUev/8nOg1fyjhNm0fcuO2k+HxuFUINQ0hBCb/cLPUYUDNEGBsVX
JQMA3SruNDdsEGSqQvgIOTKY5SM/8Y43qK0gFxHPiecKjErbvmkTJ3U2aoItXYjQ98dZ53H9I8Mg
zGu21SFIkjWM2EMt3LkR4F2ikEfRXZQxJa4BQDSe/vOD0SgLzy3yRManhASpRBf2sGBVpEVWJ7D3
EJULdOe5l7N7p+t8DpQkBt6nQwV3hBw8VBv/c/Nc5RHoYrr2WzL9WUF1J7/Jlh/nHquG9wxBYykT
w/lrM0zNZV5PxHjCISilkWnRCopo8SwVO0uVoldGFSJuzicdvEIgn2y2xiKUFq0yO4/JcfFsZKVA
Vpm4jyf7I+cujdJyLai4pEEn5ky2hi5I9ZQV58Tlqbhnf2rKNbsZkg/2VtL9rdmFpn5zEC6kr7tM
lFbLjsJTTWsnFc2iGNOE3HxPbNGAlgx0YwVbTsEnFSykoUkoIVTCkuXev/xKloxdK/KiXhsCGwWI
rC+okqGDWuiIryY9zQAS8ttQ88CMh3z7Sk6ZDpgNo+pjFyabTuD5AsO6F5Qs3DIzv9aFMkggxGKR
V8uZKolv1rMFYfct6toG69tXOWTQRjL0NRjtGZe+9t3+ean5nlej0IkKPQkAMDOwrhvlUxvO00B/
dV/knfHEtix03QlM8LR8C6cBtX3xz0ER6cl8hVTtvj+gud2LQW8H6m8hmsxuNcvCsuUvRgqbJRV9
jtRf5BkepOixMX1jdNRZHi5/sdV8j/otpB1Pieb4YeDOsT8n3eJO5EwvM1iLQI3v3X+ARgXowGL+
YpNB7IY0EQWnZ5Gu2FQIDSrNlRNzLyWtGcLQSKSZKS2l8rm05ryp94xAGtOo3nunJrL6OGTK4v6k
aTvj3wAcUjb1q8/riX7t8OiMcjy8tr/kyt3dw38Bft+K1bEHElNqDXrrFv5sz03Tm+s4ikP9dOrp
pAraNWRjs1Lh19B0l9mTtZY4Xvcpd8YLJXYw8BygrO+QN7coQ/wwSveLY/Yr3f9YnkvjXkAnwWDm
ccEt1Lr5oZEAsmurFScXhu8PSf39FeyByN7YMI3hAtQ8B8mQyorAR5qi2Ui0K0huqTtAd+cqQZl7
tOd52r+ddgga/MsbnyP3CNXWh+PCmBJ5zKedk9IbljDKsJOQqNJdwWo4bRbRKnrzbDObQerr2K3L
l99ULnJc/h1SbEtTy6SClE+MKaXbaKp9xMwF21uceG0TvEvwKi5Vuwp9qO70YVYQnKJ/eVC4stF+
21NQpRe9PKPRiemMVfikO4Rc1y0chbXJVRFuq0seRUT2L+iYkqBuz/G4sPWWLB3KJ1LguvLLM9vB
0cXZ1Zo/zNKA2p18ZFk7vTe4AkmMRgj390e5F2ml1zqGj/6lYXVcJUp7H/OXZ4j3IaA5GbuOkh7W
vLKdsyIf35HICGNqjQr4QaP8NlyFvAVbzD8H4Lg5PVRL1F25wmof/+lShViv0pSRqDl9nDyw1D3S
TzmnySOVhiB5IqMBYsLQfxd0r0qa5YHJMgkfwNr8vVsDf0AI4JHyv77pxeu4UeInHVrwb8Huvlh3
0v5NULKGw5btDSfUVV4boIVg+7ouiqxC3kBCYGSWREEnLk1zN6lmm49DuiRadI+tWDopnErkRdh4
7WTCgBDPK3vGg91htjuIjwZyHRYBSPakOun4tAqj19a1BkIZJBoGnaqCp4jwrG4eTHrlyDsgEtWb
qGZ8G2se2PB9yNAR+LcIhx1tdcTTmqTMRxDHpu3/OyEx2KHp9Z1C48kcw3SeBoAJ+qz/wPe76c3C
OdWaE0y13l09cvO4esRd8Jac9mF1xWVSyVlLoKABAQ14EHaSTfRJNyUzDFsydMr33cCw+uXvFP9g
GogURCc2ZxSMhSI4Jhj465AjoqG95oFqsycBIt5CIVEK6l9Kn9dlul6JhOONGoTndhajRfx2CPnC
4H2aNETRtSTDqLrsoDlUj3c46A70T7WyopyO8Dy8rcOIcQ+NLflZgVkxVlItjG3AFdPwAZtirYy2
gWMi5UShvgAtgsUQ5bgMu3xD4EKdi7FjThCg7MhLJQJIcJeevnbw7G6OxHQXlLeUEC6HI3LxZyhj
S+jbhlze+lD+pkNMscWKMgCLHfgoqzPX2TeFND7O0xmjteroikbqJiUrcgjMrtT84m6BLDsOcOav
qv1rAhke7zTccYQrTTdU8kCdPvYB90MPNRsLUjBfpbjyQChwDzscWcv0ZaZmpta//D7z4+OvFDDT
mlLlPbzx4QpoK6X/1st2UNAZr3+9kqGRwXV6NhRBYNwwZfwMsnb0lPxRVrLfadF38bkV4L4HUtBg
RVM1xPxLJc/R7aSTODjvqOjwO5TWR8MegC2cX+65u7cQMphYD1v+8C+Zldvxqg43NJo2MQBa1xmF
uee+tIG2YMkulxJk/tsIwoUjsxkjhosvI4fqMrHtDFpFekpa+2ONJoO6KTgsknPqsSQTXmWQMy2U
EuRTgyg9jbw4lMh5xkjvy2oyIMDeHDSTPFD17f4LIJd4/Az0Gm51FI0cSCDXZBbIcnknAd88k5iH
fUjq54Bvgc1jlnW2MyxYsmT2XjBqTfXh9UGVXUFV1KpN6m4FdlxsDdg/uCJuWFSdAPC3CX+7hep4
mkh++XK8OVuUkN95rKXKyYS7/4oBXrrIrTy9shdWc/OaE+0iNaoj7tV2FGpBcJ1oYAhvdAc17+Ai
OZuUaBG6Vd1TrPBU/BJLE88mB3mcUcNwtA3vVF1gVd56BMh21hDubULPxGHSTlpfccJNjsDchNgX
tm5gOVK3lIr/f/fqDBTM9Nm+aCkT3WlO7BlnOZPqW/u5D/4sy9aFVJdwALnYTCk2m+MqMDc1p4mL
dGzGh4uwAihfcgeBI45mUXh7HQ9ZVvhbFrcgJ+FvNl1+6xgpr/wuNV8vqJCKO+I/PRB14/WgASjY
6gcgUUlCH9ei19HnJRcc8UUp43Zzu0v8TOFTl/eVOlhWv453OnOX0wnWhzQxsIlLO0YCw2kfUxOT
tRuVH+p//U9DBfcUGiDmWN9I0HV40aKHEIIa4ItEGYWc6a5NdusG4CdFmnQdczZtX+aWkFqRsPIO
elDm+BUZy74jtTt7sarvxSu8+T4yjNr22KqeGlcOiO/TXNNzm+BeAPMSamMaDMih/EtLvP56AuGK
xcYjV7tm94hsVWr3xPYgxeIvFD4ifiroMiuOtXMlfmfbHCwB6CUPuyZYZu9RBq6rWLv06qQQSGWq
nyM25AVaz6ERb5QBmQLdf3u4NxF3RccZuoFbo2suMoaYa3y3/cNMjggxMVfA8mWPVVEQquGEVMBF
kSwE8eteLb5LXbsXZpetQDcOvDMSef1WbRPDkK8rR+p+O5JXCssRj42121E+EjApATQel0TI81VK
nGKrkEtrQRisgXtNVJnE3Tq8VQSVYKsLsaZbp3GXkA4pzeYB9gLNazkiuwI+c5hmhgI+8pP+sSL0
laZvoPA0DEsNpFtMTFIR3c56wAdC+gCYcq/CxQOnB3sHa7EEwVaQ9gMc54iNoPGLcEdCmC4FDJLO
yXkHUDlmg+cjwYk08ndqZpQ6z/c0NjXCl0mQdUWFBHmNsmQpnWp1fo1rNvM/MQsyAIUPTdVTdHv3
P0xZZz+1XBjJHD0k14k6YNrOcX3XGYI7S4bZfKslXK9xXhtwXj9yo1kqb0P0dNZUKMz0k+Z72GzN
RUj+gt2pT3PFSKJCinK8bLz91gXYhmPBhyRjN6/AA9sRJEXAkvTD3YaKi8Ij0ySjcJKAldzj2Ww1
gLiCLTZWBbdwXnbOiPfvipBw+b9bJ47l6127peanO574Lb4vgtvlOTKLLoMT+/alcbffX27lebFg
LOXNhwiNufBGLEtoMW8DduSXCEFItz99KfxqGsyYGY94PSFssgS8HvDPGaTZJPKaEjc+CrKsTDW5
GhIiqxRj0mk8ZQbck2dt8LDlgPCj1ZsfqHNpbeBIoj4Icns3OOt/pBZDf1gqC/gV+jOvWowdYyrj
1nEjN/lhx+ME7kokALMGkBWZqQFVWNRU+qpj5u1UuY+qtLWWRBoArgPiMVTK1wG4K0x/ND3FTu9q
tSjYQtsj1BQAFk+przLE395pRoaFW+/mZ0SM9XUw+UF1uPmLEFI5Lk7up6cJ9/MupPRnDDfSA0Li
ylJjLlYATDGQWWZPSoQQNA/UcQj6IEMi98DD4gd5cqYGA33SQXnoRSPzBiM40oq+P6v1JndIrD/7
7nfhf8qP1k0li7PONWXypiGi3WoGi+NnB3kZPqhqJAu1YHQGXsTwKWpsHaYvMUIAPLLreNLTMb8g
aKet0sPzshPCri75lL4uRlXQYUxRXWqqK4+fDevHyC9H3Vj5OnBQtwNfYWHE68L6bwDFTaoKTI/Z
5hr15CQGFvkXzyd3cWkeMME3VVRS54D+M5gzUo9HrRkewRTeaWNgE4Ybd5jmRfsJXUyNWaprKjRN
BrqfQQPx1PGHYvsFWJhaEtnfw3IbfSqH4+MTycjUQv2waMdLOQTKW0V3PlSnCb+0xvSG7xNVMlFi
hIopEMcysJcpf/6hl884phmvS3nhjCl2qgnPMcCT74RgkHPl8WjRT70jEfQrrFDvOLtMxXWc6uCf
9rHf02n/aESPaHEJLl6Ouc4I9g/BQflk3WSk3ro0q2K8Y/PylRTyyUJbPkJPZI7UQ7+NrgSx8E+x
zeRDxYqnSZZj/OdSLQdI+qImhhr0tOCchCTwUWFQ2y67QlkjFuneV89IK9CNqP2eZ+aQLorPk6jI
IXrZh0oGRwfYNEVylAoL5iFxrJBBV5jbpkk8n7MG0SBs3LLzZU16OFh3Fi+LN0Sm1B6aRFdhLrKV
vs+6p4d4j4AXGvinZKKd5M1ouig05KJx1zhNP0lwR9r9y/WFj8dXJV5RXjoZWMUiDpdoCwuDuOrR
toJxQxKxhKfsa4xZdKHII2dERmsxfkNsVOZctRIsSDKFoo21DZ+ArHDMQuiAlIZde4t8m0Ubp8iC
fLInkDvQmDOESl86c+vW5NUG2bxATUdR/NVfeNptIn5UK7s9X8IS2oaVR0O1piJyggGBs1uMMPeL
ZIBkmRAFf5UzrsdzcpBTCndUg3/Vg3D8IsbnoMYNaAxfsbz/gK7mJ0SvIwA2tAXRJ+Q+a3DNN9Z0
6ZoRyZhBr4XgTKAUlyRhNurj+oBjLo6R04qslogPyHrXhGnDavi2+A1ZVOW2kGCm6JxUb+cXQ8mm
Pkhr4PvUeBFD7T/KpuVZBmfaTObPQopkup/XVbG2aql+zcH4OQR/acQko6Vib7UFkeJEXUhWDgHU
E0TqhYuZx3273sSc8sgfCivvw23LPLNZBAmyUPStF2DjOzskH+sFX6Xa4k83cAt/b1tVVYuReVMI
9NpY8GPNAJsCV66/AHme3JkFYnshMq46gGoHcpgX/cFxl60itwTZ15AbteNEgHJ5QmDxJUx7cA+N
g2sIlYysJlGxipZMWdpvT3HHxA9k1pbUXrSEfZ2nn8X6gIk+Pe4P2vd8VUcrtJLgDsQ7HxxNOQc5
dk6jGloOaFkRcwdVtiBHt/jHojTLYi82i0/gl9ab8jZJpq1RVdUemdTglGmVLBLLq4ztoUq8LYLQ
h65oOOiU5pmTdAVnpPWORdlqk7+PjjSz1+cGuo6KZGrq+l1wGayCW3WvhEqvdObTAa4TYUHfHr5Z
NeTBhQXsLY8JtQJ1gwVCZGc2mtAZJSlXjkHBJFC4ecFFlF4NJaMdo0lMYXFmOcxeGuC484W8bzhr
rMsiDwfJWjXginHX4737NAIY5DKt6wkX2Jgop6bs38iiX6i2SMSpHDjiEM9Ae7IAi5WJMgvv+vUY
jKKXLL7NoHcF7hbnxVN4H87uj9DZj3u1TuyC1Pd7UKZHL5yk1WminNV6UB2U69LXhO+39OT9JXCk
Mk7tRPd9pRIi02l5wLsh93J+k3OtVMxm/VAHTk3NHiljc22fVALW2zNu1CHTZmaSx/WIyLR+BhT7
+BS99+6fkcLv+1VTOBwsAHOFybASmiE7uC4v7jVbpVsMJy+drKXlwA6Lwo+t8ZDje5RFgsBzX9Vd
+pr3dWFS2Rls8Fp94HkqhCJ67qk4Og/8SoXqnjO072qSsuY0/wknhJvvFdxx/LWYtyk+Bav8rQJs
PWvVkafF/wvyBGcmu+xA2ZDmjEsfGs/M1FMPWhkKVeMM0Fe59xHuYY4T1MARKA+57lfEuBNEloYU
i4o35gnl1+UB9J0o1Qh+xR0Tz8UXc4SofbcsY5Y4gMDXYAwld9CckLYtFjYGwHVY6YKl8S+4uBWE
ItaNDSx0ZwfY4peqmwdqQbQH6BfLvYXc6KSpKz+L1dTE4E5Hw6HiifhvvOuDCw0E+zj1uzYsbvXS
ND+xj5042sYp5Dk9Ur1lLv14d28tt70lgdVdDvd1NNA4d6Ve7B85s6R3MW/enKgu0C8R7qb1Qrdc
eXu5UsnDCZfzvveak8q+DsWvm+qqK4oA3/rfGu1+/zT15lpIUvdgfCpLnM9EifBHxGaeStoly/8J
e80HVBXqU91PIWNB5/QX4ozHZS4T07cSepizXV4bNe6W3pSjZ2J57maqM2l1vWANO7742S1klGLd
kWQrpl1UY8s4fWVwcM4oPC+iA3dEfi6l2IeJB2MKFxZZI2XEafJu38uRFLAimiJTL5Bn4ZwzlfRD
RCTT/tMgTWbOjDxRYbCoUOs0FIugGGC2copk8Kh+A3EPpbjEyW8rliHKrNT3zHJMdec4RylVTFw3
gvzwtkRT+6IcE+KLrZMbQP/ii14SF0HYX2MbDF/K/7EtZUrpKtJpojWWAWDvukmdfX8j/ytca4uR
XvWQCv7p5Zt3gzIhHqeXkIsJerRD2mLb7YUlYfIM2bIf1MLWbbHIkBOqNZousj5m5IH1rgXEYJT5
1g7ZzYA7vuwmO7ap+Vn51vfzNF7H/duaXAai/Y4fhze2S1djU0Pq87SAnjG9/8iiSmj/PGjJn1GX
bkpWyK16jlPI4ddN/1FgoZZjwaUyQ1tVXOT6LXpEdwag3Rx3Jqz81XloOrnz1B4bl92agW6TX1PH
ovPdBvtW89ouZgbZHZMSgjT+ohb1p3+PJqGltG+8W3R8whqm1/YHaXIM+brnxkKFVCfQ2MMPYv0c
r0iHdXM+rnt3lsksibe4FVQH81/yb0/p72/l9CZ8xEVU14rWgXb5FEMCcumvePLM6mJHoW8x/45f
RPTAYFEcBHypID2v/rH/2FyhtWEY8I576TLRicl1sLHtc6UNcMnWco2B4pbFplk415vR9AOK809s
86kKcm0n7RPkt5H4qD+xG/CH0Kr/gvp2I9ZETu52hsxQT59reVXJlXYsc3YH3OUL9kdc+tKvj7bL
l6rmzQJ4loaH/eroOJWKD6YGvlj1ZqmmCjlYhnsN3Tdh26Nj3OGdLTUh2BEGWy+A5DSsRKU/8Jtf
HRzaDbGjQcaABqvVkU/IUKIbIHuwZfwlL1fQCJBZB9MyLFGL/xbzoiiTwjqg9AfDcW5rnjuXGdsX
oXpJcL9e9tsfWP0g+QwE01vghWCUlS5XPy6zcmUWfAc17CRfLfTHgF3msO8xqNXhK5/VNICoCcwG
Afb9SxGsc9LIbs2QW58foF3Vl+O0uZMPUw3QTmLn36RLxqcWlanzGXSp6Awig9sFS1gGKvF3fpAm
Y8mc3dv+6JeYTafk4FKtDoN4+dBNIyNfauT35wzqfxgQfeqr2cVEAw9cWEjHXkt0apHRxNqV6Hjv
LbFYQT5uRedrEFfzGAKVyFcGGynyhxlUS7kpT7btaD+C+IOIG6+V+WNVkdq0isvxnYylIxEo1SNs
rzd2Kl4n/yxuqEu+XMc0fbQvqeuEAS2D+PwW4j9+3VdAs8D5cznWIMw/o1ZVlC+GNxQklgBehGKE
9pBYmBnM5Az/tDg9W26K91cGIzDBLZR5LY/N5xSN23dSceIQ4h219FtjlRvqLrCYTSYVuOYS0UOy
a9B6PilxEg0IaBs1KHHZWd8Bvl4QeU8kk7pk/ZDIgpQfLlIzVn6F9LnkrcWiAuqv36aUqKq6G95y
zJJY7tbnqSS4McvX4ZDbAhvtZNFhrXa8MUEZVnlzUWExxhFqx/RiTvSStYyW23TzP2fMTBjFMdZG
jQ7tsDz9x4R8OUfx+0tWNHAkYtnETbEsW35DpMOmGugEtwKP/aUUWWreKhEMOXWwRLcjginyEKwM
6V0vv8VrlXwOa2X6zFDeivoQog/vxtCCKh3DiGxXpAPBPd6Bt9hu9dz8Zw+j5Sdj3jA6BtsO/sTV
mFE5CtvF/OCj3kZXPUfP+SI3Od3PAtgh0Su+QH96n7fGdbkzzbsPKJyLOzwjtI/KlIFNq+BA+rxc
zvJ5Z4VB/nUBafbSdD7HKQsHj6hxqKBV1hXI7BdrdYEThgm6/Web8HqE6U9MuVrF4/YhQEkWPz/d
UWqrdpkIsPbr3cgFrJuWwCpXX9NxLzyy0RfdtAqRaS8BO1EGTz4YSCSMsYzD7GAPzJ3++VLnVXCR
xUTDG7pUNicqvaF1lRIuZrqcyuqSZ8k6Le6a49Rp+i1Xtrt/9W6ezOK0GalcaiXgh7TsBe4TrPn4
YF+ENuxWVY6s+J+pIV5HaCtpqmxZHr9mOaW1eWqdOjvcQY/GbE15/wLnk8uJs67ElQoBp0r4pUYD
gD0rn9NC1ZjuYYiVHqfaVUbND/FCGHwTcMf/jn4yafKJrqkhVyuJ+LB+KY/ki9gvsbOIwn8VRjDv
yv9JetkizCf9agqqeZ+Fy8OQdJGnSs0itqJ/u1gdV7t5a/wildIpGefa6IGAXqRGOnWyh11+JPDi
8jclQdYlpvlEnc8AUrxKTB37/r+Bqklwok5SxyywoHHuxwQ3OvXufXBifD3EdBcgsePXid3/dIkw
9K1mALBu0vB1IvWtvsNNQfNo/QFmIu6npaRZLWrvEsEmbqEmCTTGGSwbJFbbEhNfAAoW7TP2Y+gG
TWJdxkPDznwFGSQ3Acwp+MNuRfZYzBIMuYGylwn4tX2IgU1PEZsZD7JR9mS2WWW14JqRS5/I48BD
ocGdqOCA1U4VCaCGARveWwLyDdcJfd7ng8lCmonzx285O87jP/Xifat18a0vUPGYWxnTOHAslsCj
fAS3mmpl5VP7RDmI1lRwfS5j8ICide+bcAEAKgsPBwfE7QsKVm/0IbVrxnuZNqWV8RNXhAsqOq7q
Gssp7aGWVOjVdy0d3ilcMauNxKoA5xqe8i11AID4E0GY1edocOyCKePc8uadeJJy6aD5ZMb/Y6O1
TLUB7XE1DuGj72dqbamxzs0qHp6nTTnsCZpVkR2iK0SpcbKN5NyXKRVEpnt7a7iRuQly57CilFxd
wnflM9zMvNM32lLpQh9jw+rUxHt5sW0bpo1RbpMEZVlKPgaQznwcepcXnzrXHERpqWlz/SLVOx6O
u5yaZ1jZ9KY3JT2sFPEe396Vngn0miMhtpqyOIZSflV2ePJCEbac/PUR9b2pMq6qVqzpmcgbl4G/
UQY1XxqNNQj3fnvRgz4hz7TwEdmYpc4i8tHycwAs5Ys3DjZAywirZuVVH2bnVUCKmThFy518ACS2
G7MIrz4QzcGzuV9qQf8YCozwkHVl3Vuf1UWA2l6tdAlEdfLQgfs7fLd1ZZSMws+twfzlJHLU0P4W
PEM49rYRLDJQRt0N1mz0Xvw2HZDORwGevVclOu2Fsdd2Vjc3GTq9l1guSZXRTh0qjjt+s65LfLU2
ueqmflQfNl6eskEbscxYSbbOkBmyQcXYFzxjj16Qeoc1mzNnqG5z3jhbO1DwAezxyrBrO2d4kML3
uc/kM0DC96ILQvbfitb/0m/shpUxnEMRATugEIOKU6mAKC6xgn7PBxypOAcLuat/TPgmEtoFheLM
zMSh7Lks3Za+vxS1kbC3/t3UIlJvy9OHVK+EPsbosfi2W5CYEeV/rvxURMcrfWHYwgX5HUPf85rZ
q5V/PxGXQFC58wMolzh/02Px+gzBqQ/ADXqbua6UpcpZZu8woBL69fAGfe+E0rHzb62CSn3Y7Ssl
e+FeN0vgw0PFvD+o86MfYPVXNpDtU4dQLXwLMmVc2mMLjn8hqd2v491JQQ6XFGpyvsLIdTjGL/iG
Q4QS5vZ5OKrTeXotgzLu4KFs5824tIEKMt3l4l9zT5JT8VSwgReohlZskHIhIuJBJycQjfWWDePj
GL+LgKL3T+68cNlZhinsN4j7HtBkCdE+NTVFA8DdcXpeYIruHloE4LVlROTvpRUgF3jvZ5ITL2om
uBirhaUrnejet5i7yKDh33J0PJanq/ROGW4Zyl3wBPpjQefHEKe6btQWQ5N0v7gb2DDLXxcMKHFa
mvdLKvlEWK6+sZyb5DVO8/qjshi0zCE80pwNqy0g3wWetRw/YCFtjRc5YBTkkgbwyBlQ1jvvTyla
diTIJpKGCAvy4rQJj8XZOIFqqMzd7VlRi5bPY4kgqa9JKSOijmPf4gJfNcsjY+t83gMK+wG5YkQj
mAk4GUuK/YCUpa2dBGZeTTcUCLhJtDf1GbDR8LUYV8RwWYvPP7r+mZAwW7Qv3HdmoYIvA5U5dZfi
Bdae19kDa86hR64BgqjNrqNw8RVyy1LrijyT8bz/0aIwOhAONW50L+vg9z7ndOCxpi1TZ9Qt5v1C
e+YEkqVtYwueRLxemsk2wHv8ZlWRkJdVQc8TgfJFSDP09UmDrWSQnqaiO+H7dDgZWHJblnNJqCEu
rOO/CxAA8IUjYHHb7U0m8wzs+W8g2cLN2VicNRPGMG0iJKOtj0semPjMQ/a2LzGtRIZUSlW1S/xc
CarMBkI3nqZDpX0wIol7nqNBijgtvT8lv5kQQW7hrPWb2g5bsdp5Cvy0rvAlxppfSbTGvAWnyJ3F
DfXTMTDhoqzXhRt7gNoqiOo3P/9mQa20zhJ//XW8hmxHTQFtkIlWtuQpyXHCwit9krOGid9z5MiH
O11WBqzaCd1+vPz7+qsZQn6KOe8jplfmmQhQFrw3+/OOR0NyqrAI/PtoBjoCgbl91ev5796yCVO2
R/05M9b1fzdddRQ5lDCTVOvTBPkE/2nF+Y3YtS3JA5Fv1GkiJY10C9crmcYWzaVmJy05ZrD/zjl3
ID/ffzJSQCSqnhHQmTOf6NpYcid6tXc8ow9mK0OAYMAzGKSUy+KzzYLJ792uDe+e/D92uZY/2jVM
I60Pdx1f4pyg54OBIz5TfPI7O0QcLe5ClfR+PACtzyLNZuRx/uojQRXSo9VIUBO5BkyaIQE3973O
6ReD/Zn8+/HqufRXDlyRxJ4r0l9WFahE0cSHFgMH3nSO5OxvQuWwLf5ltv5hlkefs5rG34g62kjN
BdIAm47PVhb5KiLMq2Wtkybnp+oUwduCcfcrXhto/gfA3nlyV3SUdfjKUybr8KNsfkQGWBhlfaI7
hhOIyJlhfxfNwNxPBVGXWAe9woRqeRtXuT5oBGAhai5P8pihSeYYPKG7rjmD3UtEj0O6yFBOZduW
GlC5vapTlC7o+uHR17YznVrzaRmCJDoPpqUTH1sm7QoqKWximtNlvjfUqYKS2oD9OsGhZICTliLp
gbJc6oaC45ayrL9fIqrqD6WXkhqhziaeTpG4SIvjy3AfNMXI/iu8ZLDNqnI+EuMpyzclIJMdN+ZL
sn35Vua2O2QbEFVWeKrMXe+BEdYv8I3Wd42umHdCYtH1QZa+uNFpMW5LAmkZUGEW2EHXiVt3qcCL
Qg+DDNW49OspVo+a++px8GfIsFLIa6sIoICik45qYAdGr7JZbDnk8F8oO8cVIuHY0QDKQeL7a/7J
MAjE93r1EmfCwRlJFIT6NV3PDe3U0yyb8pk1GmvZoN2zRA6zLejFj2B/qqfyONWLhSP/DJJg9tL8
DWipUsb4zagEvphV3Q1fLLfFGNDAvwL2Fc54+7MvBJZ1SoFyaYqlbWfoV4dlEt9fW8Rw6qYRPkuh
OCke+qvelvtzTcPbK5edOcv/nIqnXBnkYBcUnBP+c3rxFQ1z045cLo7K+6o6yhAQJXr6jxS7uin9
HrmBpC66VHpO4ehQMglY5omNgiCzSkRoXpwcWlTygj54Tple6XvCpquyWJ4jI/dIj38/J/H5YWNz
zeLBT7rHG3LHttCq+8sAzCHJpi3Q/CnHOvOZ5cdBLewzcnAS72mORH33av2jFD9nz4MpXKarwZo2
xbWe+zdS5UXlVdI+GrePZhppWtCx+liN5QJ5/940/RB6xnfBFyLUP2Cu6qWWCa21ziEQKgFF4oby
ygpKWLN3hlOxnSre4NB428KKxvaBGf74LdUM+YQ1Gvn8+WtA7ZlOoBPqt5M5cmiN2S0HXansu34Z
as2moTFtQNmt3cfM4oJvF2uwUrkIQqwhgTav/cVXtpXl1/YF8f2OpQ8gxi+NKgPgIwYvVMFIlc8F
b7Px5nIemwu5wjGyx6gkNe7sJRX/irz+PermFI+mc5rNKAS0ginpx1T2wo6j/3/IXcq3ayJKKB5S
rUEAVXjYvkhLVG8bV6hd69T4PN/Xp0ST7tKv7f7mbx4MkhyIe5Ku31BaaMGj1vabb1ByimO73eZg
/lqF+x0FAuDqCl0uX2waKZTCZBmNKoNno/wmF3/ajRHhmQnMf3avTXfwZf44/GXgfqaQ8APUSU8N
xKpAOvaWFWqTZTX66fKIUFu4GhBdJkMqZzye/49ew3m8a4YnL8rnnBm6UriBDwkWebETahKZw8Ju
8AXrKPoFA4WOd7+GmfjZbMwEA/M2SOKRTsg4w92z4QHe5o372ZOHywRGZZqqHk/Q2GCCAnpM982b
QDfiDt8rVWRgc2/3jayy6zICEd9becbKhKaDDRGxXkGtZ3lO6i6i+HwCl/NkOqjfYcuaorzRIRVB
rLVGDbOOeCzWv7cR3E3lZXkN0nXSlK8nJskvmEsJJ5pJoj2q/o08SRe5lclnrM2R8FhQiga2Lpph
dFxag131KXGcoElZuayv/Ymqex+0TCbj4Ii5orbdYTqwvsG/RxE6Ig1sgcSTcgknKc4j/cPbGrB5
oNfoswrIW2Y6f0Mjn4Ir0bNNH94NRbolAs7zVT9/6GG+g8OyMsNkCR2xeJ9ntCV8yewFfNSp0XE9
FCl3WYaCfotMJ2r1kk/Gpc13YJnHjPDHQIgKc7vRF4KwcVrkZTPn9zpF0tYrwd7M0rUZ3T6P5wDn
KWw5sGsn3/9QRqfqCfL2Z7uaEkDr/qJLCUes2s3EKLvOxYWv5j3MNfz6iPEl05NtNWLiw+9sepmH
r4pj0LlFSwaiijGw2lMlgr0HGXX/pA99koOeJ8k9Hzc1hcPVudDQplUrpu2WnmaL9DdFnr0Irh5n
r0Zw/HrTwWVdBatoMBEwxgOqrx1RoPBah+qEDj1719U2i3LM6uvJ9wQeWWlAJ0TLMx6yh+UDww1p
ic71aqWtR2+fZ4XE6qQPSYPhrzxcGVQfJhpPJE4JI7uAK4/pfRPA/ymYhGB93ci1hG7BX2Vwa+Np
/ORYuEs+ozlZw0V0SSwqHpVf62EJSJxe/yYwXsPibJd76RPGpgHEB5ze6mhHpti9pouAgrZeeZ9C
EZo0WRbZdkLJHxCoBnqjaM8WeVnElYj9CCRlxTP5D2PMu9Rol9wrR7Ka8o4Fchuqlkb+KuKoXEZ7
s9PljYEhTqVoCFskexB/JIvYJS8LdYzop8YjEr2kCyovLWD3ZWR4VlsFXotb75J+qNG4MUNAGyP+
OWHorf7H/s1sFMD4QvEwYnaH2UFv7kROuoMeLk2UVlSjNyKZ25kpwa0py41gnzVo3X4GV7jTdgfm
ZTvspLiIJU/w+mDdhT6p+CClllpmzRGCto9+F5TqRunMcpQmR18jFZdzDG7nfb3rPyIfWmqmeon0
SLrTAjCq3+UPWl+y5WYTgWAVm+UecwzedsH2BugyK6e6XQQdrZUkLsGM+zswq606VNAe7apPzgyR
1InjZw6c/7PkzYtFgfRF23Hl0so7Af+rWBVyxiQYEW2F0+e0X1OuLxR1BLiBUI07iZOBMuEqztgI
57z38tLHuT2B1euGPKep4i4nlKyfkUz1t1u18SzPZQy7bosAspiGNITUAISh0HcqgJpgS5f2t/DF
27lGf2wyGiPjcQevFTDEShKiwODCoBOYCZmdMnilDrjcc+E5oraDlG+ifuMClf02GGbohIU8jKBo
PQuuYWcpwQY+LuulEwFGv0/dKD6xOFnjY1fBZdYVUrXpqGbvqC0Stxsg3QyAvySHLwzktWTizk+r
UgUjDFOqktqEpbsmDeBKowpw7G/nj2AiKMLB1Dq+pu7GWzSAaYyMzt3+FTT2HtbOFsZAd4b5Bft0
iimQjYk6tif+7ZEHOD/I7g25AruRuZk3FvoDg+wFLPyxVaigWCQTNhleuw72QP1Tdwjz60U4OxaJ
EwSZaBUKMKsxK4bpaOINPEw3LQ5A10QlbhzIUXdKVvF6veqY4lXlk4vScslInRmhbFmr3X5p3+8r
9vMAqbEBLoDYIlIceNlaOGcumxYzXvwrhrJPOLY0TQjlIO9ipRCqwYkcpORHjbxWOHBBwTsbGdjK
kD/bUKrfwoWuQG8O4kWvlD3Ptc5CQIOEwWeBZ40+y8Fotc1SWWbhwVQ3sLQvRHFaNFJN7PDRv4og
6c3hgRzB8FzQgJ14cGutQNZ6Tt0p8GG2R6GwR6gq/jPM9rQr11aHsSqp3VHKshvnpGOECCxZm3Ss
EALcvfy4cpyQEO52CyquXfCQ/unykAhh5G+VGQyvKnGpK6cnaZvaW2zmNXoxokdl1TNfcpJMsE8s
g+nppgTxtIk43I6QDGSrZThiTunA07aKy26jmSHTj3DbJ1hPfB1QlQo9gJdYPTX6UXDbGwm4yVcB
2lowCxXfMfTiq3u6a4U8vmKoPW20EQEXpaSa0t2QQeaH+BzDi779VByAZ5N/nL954qsw7N90/dkJ
QgeYrZ+WooSE6+4f/zMX3oO3OsHsa+Grvmqq893x4GdtJHaZ7X6CmoBkcBU/uu1gB2pZHcabmqGx
rIvmRjZRABDbQdDTq7t5wDEZgbunptQWbn0OK15M8RwM50gG3/LVynVsh7N45L5ht82y/Cm3a6Mp
L9+j3yuWCADM2gIcKB0zKc/P6Z3AW6NMw1uTPldzQKrdFOlms4u8kH935hUhoBKbyqNsLdL9Sd5Y
TRcxSV34IJNmFIisezGaW90pPBe2N+MjLb3Z1ep9kIuhWLHp20jT5wpOXp8i1uPejwTTyyJqIb7Y
svuPsh88m/fGaVvwZB89XuiRKEFwqZV4v+Me10Vx5MK0bdHuRFxII988Pf+gdctAlTKtbpGE0sQx
9w0ZPfX67YRj8oIsHznrGNFQO2B4ZGRn2JAOZynXBS+GdNYQSjawpLcVCHYhtESDQkGzH5AaoezV
ld3PWzZAyeIByI3osL529ToXUyg8G1B69XLknjIqk3Mm0GO5TrftKLLMr6HlVmKGvsFeM27kSgQ/
r6r7HRl4eEHn6RnmzcbYJM6Mxr2DAwZccYFgu1AftjkkUw/Awwup26FaTPB58SlbGC7nZuFOjqFj
LxUS9fbqyix2bciKZDnJWSGkOnl9rNR9Ac6eSMGZ2jJePPWC5AJ+iJp3VyQchzfp3gfp84Fq6GlA
FHhxkfs9KAmoK0shVBJnjGwzSpDjhyVX9euGshk9VHU32cjnJQN3UoMIJ19nWuFHR7mIytreZ60s
isb++2IInThpkmqQvq5AM/iujI+YnZEF4L43s4AUSE+k2tUGfm6DTqxbsjES/ZSyMVnSENu2LyHV
IbYOxHPos1JpEW6z3wLgFD137vItaF9i139K6TecHn76P3DF7oX4Mmq07j5w2wRYWaQwpeqH5Uzb
WiK4MVAH7jCTB4eA/Br/XIjamWNyGVQGkKvufzQnhQ+jvhwUl1vYLpdtkS91my/u7tF4gX5TN50K
OLEMgCPwUIaFCTpQXwl9UhA8cFOcRyhvGrmaCCVPCkXmQz4wc+nsVReOXunZe+2OnDHu99gPy02q
5nI2dHA7l3biMFL4xeMzeLQWC/wZl+BWE8OmggdxcYJZP+I1MRzSGpQ8UzTRDvKARheN6bG93R6E
NeYotqR5OJ9pDXypjLyRrRAW0hZhrOLwooIwHvyKWppoW3sIbj6HpPBq3nRsJN3DAfS6cVlc2XTl
Dx25HALh3TmXx3zAGaLb9fxmniyne4nvne06oJyjU90wJPQs2wAjq9GG2A8TazHU2qIJ0O416SI3
DwvU6Y6BXhAv6fKdkTkcxFO241U/REzdjGf/JJCjfiHocwBfWAB6NJcVXsDF0xmTAY/+TiLroxwE
HxXbPMy5Xytx/bAgig8LktEaFn435RPD+u1D98r6WS5X97ocWAjb1oqYadtJHsjQsgfLbap32kZ0
GT5XZjxjMgPiMdXP8L202XCWTjR0xmUpD9BguSOvfH43xId6ixOz0bxmfGhWNlom/4Lpe+WH6VO8
RaAE92kOUH0Lftj82kovqh4SnXw9yA8U6Ec3kUYkW0NAu9ms7oJZd2SW3swLglho5ZimkB9m6qh0
iMtTGNwqgS5U+uRlCwj5wlzwwIYELdp/SK3Bdx+8luCj8PByT14ejbjx2EWFz8XV5X4B0YOSxpU1
Op6SP2XGIS6HzCLnkRpkbG7MLLh4Zv4W8u7K6ci0ja0NOhSX+SOp2hQQg7nn1Eg/1H6Vx1jXovKN
mGFtBYtZkEjRV2IvMRd3V9/oDjMRUQ6viD0THztts8FZ0Btz0aEoBIXxUUTzd0RI/vgFUzCgJFW7
XGhhOHpj0ChIwLseWZubZW5A/TxtKQGamKjo0LxBjHwW+WvIWjYfnSDyzi4yUdXizwEwFY3X+FMx
zEXMP7aKnppDyGzVPozUg4rPitwMxy5XqxHsaBqdgWgBlCHEaU8RleZI6mmOHy/rfiRFbDpn5Qkc
FYAXE3vFlc3CSzFx5+BvhOM6dBEEoZobhOVE/sIimier8PCsoRIP+93BkTmyHAaRrVdRAKAtuppR
dRR4bJS82nakGcbDUjCIbVTf9D2dSsbc3gSmb6ax0kM3v7ImG9UrXwJZw/Xj2xhKWJgsj8KHglzd
qH/UTW49YYvNhx+lDGtUKuTBCMbALlHUednwPK+0oJ8TRBGvF3kuD3M6CGbp3EoAKeMNPbXFD1KU
B5Bb42pTMMe7Nh8LuQD05bSTi7eKbcTIUxm+l8SwI8d97UzKcE+lX16BFZYUEaZOtFFnoc4QAtEA
5fCx6/q87sZTVsmiE0IasMhcTaFaKGwTk8K64j0Shb1ONXkTwCQVCyO+JD519ceJq1hrtNCEenn3
xgS/ihBz2MQ4myt43wF9PAUjiNmOAjCePzJqpwCo5EZlvqoqyBSdA8ymyYkhYy7wVXMuUultWos5
jb7MwYMCtLQ0mLbtHb204C0x9j9WZTXeaXI61vlOKP4CHOphHOAW0JbEVCw2AcbpxAUz7ZE9ljFi
cCGL9sL59xAectxxAWw/7bo0nO3DCXX96DkG5B4BBxWZoa3DW3SAIEAyzzaXa1TanpHkZn/TFkEP
+zx78U3oy2p60YYAs6v1szFsR0qqB8Tx+BSqaICeoaWwLAfGYiyedyd6pI1w4xH39B0fjcmJfn8b
z8Ilj4GLIiYJDYODL0RoPjx2fkwOn2x3UphHBlSF5og/2DVjO6Bk5IMfa7tSnotKoH0QiLI0Y2Af
GSaOy0hFYqHpd14EfVe/ZEEt0G4A8VfKfBp30rurfeUwZCIoPi4NYFIgM88DKY1C5EWwbfgLqcHP
ntf/byH5k8/MSdkvrube9E6jhk7XWpIvERbZaFpX/96xWkgwZuJjQVA8UJVJPpAkOMJyLjjMDUez
6xSL0RNvEfhT47DXrs/GRN+FudxurJsqM4NWb8XHstxo831IL8WEYKemkw510nhDBDByglsbgztK
68rGB8mq1oxF4XTTAy8tmCVhknQUM4oa9KfuivP2IscPvtN39FGiO1lybAoc59uqG0Xx/yxMlrx7
CFVkKDm88Z+oGzx2Gs/7iCzqtj/syomWqxTWYvQIt4vfMsm41lMbBIlEAQ9KJzT6vzRW+YRVtXcC
e3Q0O5/mn4vLjGfceBVKa/3b8zGXUbGdoIFCCNkKSciUVWV4cri6xV8zCd1i8Qxt1mbgWI593KSz
BTAnQsgmCUXjrLDEOePdlOmf8xwXvQoY3V+p0tiammHp0KAlgnvK6H8aCCg5Teoj+FNjs8N901jx
P1u7fRvabUpGvq7rsvVQaWtZbXDnc2llPFNKRSoRfr5xVmoe+y+Q7iHmdjNxMqL3JYgWAUe1nili
9e3Hvp2gzJQh83Qic6fXcenGLOxC6l5mVy0SfVz/f5LV3cq/GsEons3qzuIoNue8kPupdBALdvZV
uN244AXuCNLZyiEM8DjTUkr9bkueryHiHoVcmCPUN6G+LgVmzWDgDJO25ccZy0TCO3PPruHbAt+W
cuCERzxnK9CddBc0Sd4kokFGrrG2vmFNde/Pb+ohIhQ8EbTwQbzKm1HyJvuY2j7YLZqrXFcsEuud
qeZXSwCNNIpmQP2KOJ7/32AdBenUJGUsJDZLk68GPsCwORGRn5LpKOKMRwS85/QzVSIAN5EEvsGL
98UiWJaRL7GDeIAbtygNRpQ5UV/xZQ5eYwSvjoBMeGvXT26EmLMUXIHuvYqxg2n6LOSPUhD3eIPl
LmMvDE99xzxHmmGNRDP/ZEdJu49pWjf+Ci/e9eYx4l//nszlCnFG+PKux9KmZjeYYBSBBxkviAHg
YCaeazvbga48O+LoLt183TR+lK6Afq/gTHr+AvJVU2N1zTs27gyY6LOkiTdCEr2txwiJjbprRtxq
LgL5TZnzDayWJyC0L8NKPLefeE4ZIyiNBtvxvyiBuZSq8yX2fYHPGIn1aqE264WPH8nqZoe26d8j
YqLkE5vba0MYW5OiRUN/YaZhg98m33GOBDgTlWhYf8W0eYf/U1Ef9WmEwNT76SyEQHRHXdogS97D
yJSZGy50hlgCb2JxkZ+u9p9+GRwIeqnhWRsVLN50ZJUh6EPtgrL4Y2x7gSsxyUSCjTwMwfYNHnuY
SIl41PT/dlg+mD/bktskeGU/FuiSSRKBWnl17tBcpAD+WVv8ROnZx19w54UrtXqVkpUsGtlEMnwv
4kpQKVLK/vbY1RqVppzIapx403xzTQVMk3BB22IBUZavnVvNbZvD2GypELh75WQQGYkUb5dCZenl
+aNEoerRzPrv5F3iNdptIaFbOtI7LHgxzLQAKurkwVMpqBgsXziDrEXXFRQYFXfFVj3WwwI4jSMO
xL7NuIhyJCBME7NH3zglcZeNERDR3z5ptFWSFFE04VxBIxpMZuUrSyC1ORP4MHIYrdAyfDg0Z04D
xN7xAiTVaVG/Ey/bpVhrRgF1rdj/VhowsAGo9767nIgcyXTbMG+lsg7YB8D22yGSDNTuhrsv4b37
FTeL3//fhHWGU1gxcWBJEqoIFUxmNJopnHPIObjU6hxy5TcSzBWYBZPr28CNmNNFwUJx5nWICrb0
g3y4XOH2x4jzn7r+xr7TPQlIw1XDWHSY9NnjygtYzknJEpIWd9vZOZdgfyvVWYvB1LcLxZv2/PVd
eg5Cbi//TY+q73MfD+AOEkjFOWpPVcsnbKXGK7EkYDqsrB9IIMPvOICumS/dOAn3haMBiN4yycLt
NChqfBdGqerTITf0cG3g9dvKvqnUMDNqHcnfpZj3DnM+/XSm7kMRt30uQvkfweFdnsA5wbAw3GoS
qs0NDp5kgmas7qRc97toRn81xtySRaSf+GE08J3zVtvPbbrjij6QJLrOKR9vdYDNd2E0nwmZBBJB
nsTSgb0vI9p5I7uudaSFxQAfRLEqCHxkyJTOH5NE0kHJMiLLHvtYiZDZyN2k9XOd3ropvNLqxk/q
ZhUNXUvHO6IiGbP4K38ZdQV+HPpVPCjV5jCp/FbNpL1c/OBBzJN2usA82fNcydTRCD0vvjaF/v/a
9qeVnnSk44o6pl3WNNr3zIHfBLQ2ANe9zRR23noFHoO1Ixr6ewjsj99H0nuV+nR3s1kvLwA7NgNi
pgEU439MYIpqe+7kzcieBEItqAznv1fyduOT9zpdpEFG6lGKmzwsTkszpjWxEY3F8E27Qv5UZEAz
wEqvdNPljm2UUP2CCAQ6r1heGsWYwZYtEpmwuuxN+QDX72SevRfCBiOF7bzs/U7LIh/+Ck78UTOX
7ixo+/KzrxChwGVxbp8C5q/VYkdY3DKPQWw9/TsxiTmSzFzektXCMAkLqWcpNnXppAorhCMaLi1g
5AA9GlikLWdXLkWtA1Nb6jrOSKeKhZ1VvY8qXibhG/y3dBzAhvcfoAE0UIQNEzbQHibS/QcAPHbw
BGJWX32zYc0XIG0ZcAiXXt3UDp2GoPIZTaAoEQj0oK3yFyvW5zrqyTY+v2chgx0u10060VK+KmxH
K+JbhTZPyKMcynXUdBP6QoK5n6tuXL15RjHHXyrOBe1BDH5jB008XbWRqUjf6xocVnorz8o3WxYe
pluvxr2/uyQ4hwS0JUH+fc+716CMRyxlMLO6+qkN66M/McWOFYKZiR1X7d7StiC0xoROxu+awb/S
tbXIGPpPKVTBfdKxHxeOJgIwXjoUtMjGwv/7ODGtn+HFrfX3IgG7ZmGeijp2WxFSUeQt8U53zbY/
ifoYCFCTRESBl1JlF5Z6iPBZwcHw1cgPcXyTnZDBiwLoCDMf7gSKD64bBvyt9rImPfB1yWnf8cRo
J3HXMd/Bw98DZ8A4hbWhoWpALyIqRxOsniJIk37Y4qR3Tb3RfoXo6dVaxY21QvnbPeh5yLSfD7W3
1ykauzultE6rMXe+FbB0SR3yODHXhmtNxsvPBVc7IpQq1+womzz9uqLzsr+ahTXDlmW2yjuEO2xP
D5a3UUZuHQuPjZQeQq+V/F+wgZp3U9H0D+VFweWmWm4yFsUrnvrnqSLT4ckQmQFC/ePYMTfihxhj
C0CyvBB4VZl4TNyPRMqG1UATWNOSrhf68NzjgCD0cfiEI9ndkvPrPBRhLsiMZXpr9fAwRu1tO/2U
zSjui9G29uEjxoFnjLYCQptYNzauYCPhHybf7iATcWNwS3KK2o7M4VBaMVMNVoeKH1EhjcLtQLXc
OqhBePBny4ehajuqshlGxK1U29dDnM2NVoo5BnL+Auq9BDMaBv5Si7mI9YNtP+f5fcUwuzyzEJ5z
uO4k4UMBO1bXWhZCArwMUzWEIo13UAwyDN8ijmA9XFoCrFh/r49a2agQf5SzM3uVAFj3RrPaiVaT
I3KkDNGaa8xRxRnalbtgCiSM2TGczXHlCJOUvXh++l2TTjjksjCz1AoinjBnVSBRm4wjBZzrw380
pkM86oVQpjuOngXbPDrZRjaCni5Yq8dT4Q8OfzWOKtVuNVlHSDokxqlpbLj7FztuJ6As+WsHghXl
5fVx72nh55HyVxDuSp/wmOwWv6CK0wT5gtZMd3hG/MP1Ro5ueTcZvtQkjCp+fmchi6E0BQ+s34I4
QyOpd8oVJDFkwWlw4uJ49gefvTQEL2vv7S/RTiQAriASArnoJ+TSWv/CRR7aWZJ/u0DTU+t6W4H0
DUTe522zvoVxy0KQsLatSVJgcufqDsazBc+Gwu9/jSYlh5GpppXdOBsS/0aIEoB22xI79ZsUGC6v
bhMWdZCD74qwMbT29HQvjlmeGeDJO/qAEWEX+/RVMYAErdahuWm9vNOXngnZjfQl6XIl+APmEjtJ
WyzjVNMNxypGXHPonF4QQ3kjuZnWgXWVPVzZsvmZk/HTOFyUt20TLNpb9FnYbATSrxpTJlXhoXnp
t84TizMPLFLK8I2SG8/4d2/ENyBQ2FGGb49gmZPpr2QAOji5J4r6Dvyk9c6ak/ObsbvYjsV2XtZu
zIbn8IEW+293ZvRrsu3f+OTnlfCxNMbH/ZP6BEwKfX3Uym9BjPbP4j3/6tY6mhqQW8aBSd4vtwTg
rNH+zFrA37FVaNkfy+GXLcbBHwCoULRZVw7ogYeTQS4hzSPV1DDfW0N99TmmHyYh7kWxZEnGOzK5
KDIS0hUR3d0mfVKCmmmu1bG362vtQX1fWi2S7/fEwzwEeA8KnWLAjEWgpyd78FRpwYc3VvucvpTV
QlxePfWhUmdQ/Rc3ub//i4FSO+b2S5wG8cUCCefwbFxcyf7vs1sa9+R4+ILzz1QAvFBb7tz6P0oU
Q/1aHgSgTcgPLwAAVUQlBFy2XZl2+M5rzf+F+t95Gb+6HIj2xzZ3e/4T184onvfD1FWw8Sad5VJJ
d/3o9hkIlaS43PwRcFBmgwMwBsBVq5gS4M34euWMoPjRAaBQQ3YQCJ6SEhPgklBzFkICul6H1KdW
oNw9i+RS2fk0kPYjGHLsY8ELNDSWhsln9X7HaFm+FSQKFCMDE1Z524AydWXm1SGN+ERGNd0GORE2
lkFkw/fHYeBQ+b01WhmcVGZcQbvIQDnmVICxBo3mwEsriD3YFYkvvIUTgexT0VnquxX4sPnWD+Ve
YYh1ODzaGhe2+um3msmS1vBVZ2ZlhA2MMHclj6ndB2djOcSU7SEGKGi6QNeU4fn492e87rnlDf0T
9ucOnt+JrQKhjFMIOvckPORDL/6JYfLtPFtK6keb6BdBDEzQYGf2yRiHNSu8cLFwN7vuKM7M2TxH
K4G4D1hiAByA26Gwc30g00vu7uj5/ZD/XEhHLEAyp9vkO+K15F5B/0d355Dd1gzizQZwUBJ2hBoq
LA3kvmGE+E39m7VeAAhnHV2IMxQG3sGkeIwGRTVETCowr5uJaAxbNgbahRxuxUjw53BQpVz77mME
rgip+cmpkoRx8b0EBxdJRM9AJCs0WbJUtuIWty1dJhmuvxNbFLuWq0cEoZH2+raX4KE1AKrGLs/4
o6iks0vu5qXmClkZ3rSDonF2sS8BRUkEm9k/pY6HgW0WCTM0AQXMihsH2KectWi5OI9bTMOERqVk
pBO7BdfTaOjUR0J05tWSVeZ1bQXLSHFUe8KjqVAFblUVOZE6K/Oq5eU0wqChM/1T0tu9KpfoqW+C
vj9cam2VvSnVV153/JP+WlSrWNv5aG2eqAVTCIorQcqCwgYVQBwCZB8Ji9wNYiK/98rYpZjkWrK4
IIGrPUJPub+4l3ePaflH5M03Prj9rs6mo/4cv9rEctvWt94+FTAU2G7vKJjnvsBVmf0jkdEAhibF
PXLoph+/uIjcTfHD5QY1pMCcu34RCh0r9OkJ0i21M2ND4tuPlyz+Lh7UEsDJzujR6Hm9EWtGAzam
GGs7UTd0tdIE3elpCy8Q1AIdDMAtKBf471G01Vebt/x7AVlz8UAZSHWv4fho/zKew5zanw6P9DIn
YfjX82TVP+8im5+uUaJH1LJgzT4ZYyWA+7LMCf6aH0iJzy2ERQ6GH8RsZtzA1JU2rRP2Vk+hpkjo
YOk8udZDxDtbljoTNg54Xdo44+b6xAlI2ju9oc2jZ9bJ6gk4PGOS2dC5dBtZO2hJudaxnz2IuivU
/Pq4aFioAXfG1b/eVt+CJphob85ftyV09zKZV2qDaU0edSZe7Wex4olLpQZMDLUIlmlCZw7gTS2f
ezl5RI7ALfsveMTSTazuDRCbaos8BqyDSCZSAtRgPhkGgT3ZFLRcjMEotg3bdDsmtosLGb/hbDEH
B5Pkb1VnBI0UxTLink5WDqsqQs1tkd0HQfWI9Gfd0B9hnZeRq9U6snnZ+TBI808UAIJcT63jbi3B
I0bZQ4akEZFoDlyzsRasK2FeNWGF1GeCZMX987SGPCoe8tjsWwNHPXUOEs/dVFM2cz00aNN2Vhb9
Xa5cQxAjb5hXsOJYGIf95COUX3B1HeeaN+b3/Vi6qMXGT2PHRmp/FsqlSNiBv7PvjyHTS7h2iwDP
Z/glb6qkjyMsW9m3RipuOkNBLfOHt+lbK29yEJw7tw+pjb3ep7btucdlesJVdj4JqVIrje2pQONI
DKzmC3ZoB9kUR9B1SXMxy7w6ms9fCwXd5fUfKAzDgORJeoXmGmpQodSc8+0XEBZqFm+WJlOL2ZDb
AFihMxScHuOHX54ZdCBKndF+PUlelWkRmO8p5qgxaSIFEinSU1Zmvu9e09axr0adtkcSWDv+eFu2
ISromqM6GI4aepws4f01X4PqGwyJr4n7btaxGxh2NDHOwsdofkpWH2H1LR469ijnbUFe7+OrBir0
xqnsQ03+V7zft07qxFdjnQIQbsv3Lskj1f2j82D4VBdVDQlVk5/vYlv3BIRsBkvUJC4nkWJHnU/l
w+qJWxmfqX5ZIwudKhhOCqJdQXw2ft2rXIsaeryC3Zh6HqnqESvQ+3NZzRFXBoo3s0bk4eqvx+SV
91EMwq2Mf8vuUeV9D68LPx2w9UOWE1o5hNNy49pXK75yWdh4WwxSlSM66d6rJ8rk/hpQz4DpI+qg
QdwbAQc7m0/lOd4wHP5WJs/V0zY8mRXgjy8gZmf8CdY1ZOwmQqtlIwwPqdKK66K8G5cJFblJDemq
qbQK4+eLbhrMyhlPIBQHJLoSUcXYQ14cGrIEWjMODApjGHe4SF2k6TNMhvTe5fy6STRSPDCCcmMe
VQ8I+lLE6i48NrEfH6nUbxNi7F6wmpp3TS3kzIg86khTNLFcsVugWEU0foDrAPA1VvCsQNvr1tLB
rXEhiHyku/qVlGj70/HoXk0wgk0k80b4+cgYEyzsro0G88xvqFH9daUBM5u/VeFw/hsPb/1g1YND
unKtdMBTkL//lYCbf62GGkdFSyYyL8sJ2R74OqmXr8P5Ijk9jBfVdnnPHyEqpY8ybQyv6RNwre1A
35+qPzR1Seku2TsO8OyjtSp8o0HTc8PIBYbLF4EkNSu3Ue2ZptQJEayqfQTV1GQm7/g/64sbnXDq
X1XLsLSzsfIHv2FwMgI0RXpZ5GIET8qdP72cLY+yvHg3PRmWB5SORgQ/Mlb1k5nmkhFN6XttNnHV
YA+X2YMrv8R0mOZx55DqeNqqYuWXufgMluPtn33wKWRwsnrnByaRWlSJB/wIUAHm9VstZEP6QfQf
j4CHgELYi72Iri9ulPUjy2GG5wM+HJZ/Zs0ytG3kFy2M545jfmA6Eqmxgx0LcxxMD6tNTklU4+5A
V5BjmnHaLqqRup/YGJ34IhizLj4vMK6lT0D9nNwU0DYW3+HbGefDBjNlInACv/bCFdj95/W20sMJ
QUJz/Zt2NjeN4wy3qQywJjaVTLMtpYjo+8aNWVAGB/Zfg2LjPxbRKjGdi8subbh3X9EYpWUMzAvg
e3o124UdHDwDNsabhZs7V/GX2DviUkQS3SWhiMVKZY2nLbhQR050TswNqm2iJKDbuiZO8dMbbDEk
NkLXJYhmTiL7wZ+P4UdR6XJ2lCmRdaIUvvSrqDVnSU+fJhnPWY09qqHG6p0R/kQGl/FC5flEXAe4
ztCbv0hWyxY/BaJ/nbR6Ks5QQuVxTA8niowbQbuxYWhnze2dJ+CKNLJ8SM1YMpCJDxbrUXTWwGMG
jwwx2ivLkTu0tbJ+k6CtCbhKTirwxopz3BoVUpI7zHMBWhOjbqPWsN9LSPhhRDKPLUlCc3PoX+vb
04w9Fov8SfguT7NbIvy5i/7NHdk8UhxSmzmwotpnuJfjIIPyojgm+viqYfX4yC6gjQne8+sIcIsC
AO3i2kYQMGuCSWIdxzlVhB5gnxnYRAQn/si1DozijvqioyNFrzMeX8HIGSa/dqS9ADW1/iaNF1nO
sdP3VEiEQ3u9tQRa1yR8r+Bgv1pKq/3pHVT0WFAKtNgsZAXCrBZKkJG2C51QSG74StaV4vguQ0iB
3aAoThzguLH0sxVq2aSrkfpZqijy1YmC3znmJG4xT5x88U+psWZdqpbqkBy5soy62Vkwskg/YkuY
kHdtfQ2xSxGGY9m9/hCShqQ2rIr1O8Nt4YxC1ZPVJKQ6DynQgGEsRA0QphfnpZ6H1a0BQPCGoJod
Rq+vOrfFq6tayvbAeUS7r+kyW3yaoiyuImhjfNBufOUIL89fjg82pubwtbrUxItlbQfG2h4N9UoB
KOY0NTYge/3Oua0pNnN0HxoYsxnU/Ei2nFBbzzCZwl0YRpqQWWkL9CaVDVGCD+GNYq9+1ITKdASg
tBgiJHlwOzo/CMZYlhOpyj8S/nIhLelRtGVVX2aeCfD8qykqkP/G4yKkU3s8PmRXS8UA/yFtenOm
9v9R/D8CkijlHoo+ta5HbjpcVeO69QJZHLSAbiYD6xLvGNv03mFnZgVspfswL5YoUgopm8cSc3lP
eBqEUOe11mgVifr+UrXaFvEpTOwb/nfsbb1HtrAVX4bTEy1ukNJEHm2YfOkd8UbyWJ86QoxL52kd
+iR0PsdzYAD6DNxEVfiFCl5NOt9OMkt5dRKleJjxJvUn8OS7bvBvltxEn3XRSPiEbjKMV9bD0EE5
btvIZ7G1DQlFeyGoCoQ+VjaywszdMIzI1GqABeCG+N5v2Eeha1rWT4y2afdt2fD6S4CB7zat8cPF
hNQyDAWeBx79UqTlSqkoivLA7hWzuWBfEscU8EBjGfu16EdXlxxcT7T2x9hlfEJazix0ymcBULRe
Sb76iTAwvYPTSUv9yvakhv+KfjdYXqUsvRWVvGDzTpfcgbjQSHxtAOmAlRcdIuK3tOfqpmnEr25Q
4GRzdEsJ1QxbUE39g7mreWVzN/Alg9df7ss8EgbZ44oR/Q/4jf2V2Eo44t7cDHwtZ64aiR8DZ/Pu
wit05DjYNtTM9aXhi1LEgN2C3iL/daUwsHJbStUlyHkzqS2fQ1H16ADAasrhhzaxciIIa/+j2fIr
AQkuV1jB7Xb5uHKaV+2Oqf4roUQuoS5zVetX/Co2IriTKJe6d+qnTrI9qBLkbUNGEVitwBEkCTd2
MqutyEpbq/SrNS+WsqnEj6tb903UwiC+SurQ/cisHZsjuVhojwnw46zaozuPBiit2taDJqvuotLl
c1S9L/sTOLmthWQeE7v+BQcaD+EWFGXrt8FLYgQ841WohSHAq1iyBWdG5JnaiRU30tIkAk8lP4mA
Yem+EgK2BxmsHo8CXTcsIgt5OFSmCol5wJac0E7coFRsjDEnyMK6Lnx/LCuX/eECdn+Q25r3B7Ba
O/WfeIsKL8LU1CqpCT5rjgikXJ31vkCRQTv428sQzbDhC4lapaXA2iP1C9Vh0sDu9lQ5/UnFUN5u
eDGP/PMr6Tvqrs4iCBJ/xyboffLeqPvKPqe+7hAadCohfulQnfMkY1iez4MyXjyfKmk2mVojZrqC
fHvKymZ7poIFxihiZPdtMrxARWKeUVbdfGkIK0A3fdSbVInXLjE8Feq6nylBugoQM85mUzif7drY
kp6DfznUlRPdcKhuzgdzzHr8GENukK1K0Rdi8+9DnnBoZkxL1buw7V7hUESeVSPiLDW+V8lSZs/P
Gi0qqhOfal5oPOgFpmI1mmKt/OaVjcbWdkkEoM+W2Kq4u0/UbwDxWeQF+W5N7cubHdGt9IZ5kPPW
39xU2YOcR4VjS891WwJRXx5HcvNCmdjO4NXAIov2wxxeSeIBaktfpUJ/GNW/TN0rOnI71rwwY87f
9QixXp8oToDbRzKIvBN5L69M9YESgZMaDwSD4OmcN53Mo2xbcYKA7GYjqMAbXSXEdUmykgclfy8y
MTh1cI2lbVCYL0kS0X99wbmDo6whFbSABNVD14FuNiMRSLm5oiCy20bBiOSsXe7ifLFIjDwsDUEC
Xt+YhiRzuRi5CPJP5VA6KJqWNQjQwgK86GnJEuqj2KOeqkHexPjUdvBZTaWVlLN8OPWR3P3XE/tR
crXyvU323iNFXz2TP4XgksJJ+oF6BjbZ4s+2IoXlCzXBjBc4Qcu0sy/Gi5t0rqgX8VYugHo3A2rB
937rlwju/ZE7+44k6Ip5DSxYu+k05resbBHsk9sZ+A/uSjkg1IEKf5j3swv//iwRTIBuNCl8PmsR
qf9/6oW2A3d693K8v/Cf0rIdAk2Ow989mf1P01F18xucIUJRtCa/omHLlXVXPe1VULSncH/I55NM
LWGQJESjVfIsPaunJjG5vq+GlLnSMyxHOwBVw5RDBwuf3Y/bnrsJ0R2+8DcQLc6gkf4ojljoocHG
oHZgspzpdVx5cs7kihXZdXgHXhbKk0Db0PIc+uHi5OiENZmAIH2u2a9n80n86WG+FXMiCV2IqKM6
vJstRaAabb6y/rb8rYkId7AucA42J4ka3PpEGkRqiZ5gf8H84u5jpWQ3sVWO0Ea6rk1DMPpte9eL
obDNVpQRjc+KO0nfbwK+ZfBjZnC5Ue65zS3CYHU29EzSJtiZCljfU89+tBe49QaxxzF7s10FLL7M
luXAKQIbAJaVjCBYhj+tAykKTdAPhsRhknnX2mye+sPQHwEZU0KUDm4GuE6G3dpMAfGcxD9xuVSF
owyn/+LojLNLpVm5kgqxm+1ArI7fz1rLrFxBldJuOOZhb3lcolU7KNq36r2xdtATtv0uscvfg7yY
47tToxWxOA2xgm7nFJYOVoKQ+CAVPhNNOH6DS5pdZf/3IxOS5WhhlabobG7m3LItUmfDgIVNzUPa
GX/Mpoz0j21RTMYKbVO0CxaMx/pz9XRiTbV3h0XtC7JiWHA0ys8sIonQddN9tmSHAylV9eilCe/u
Hn80pcITqKcqm/HvXle5O7DEvpQa7xDfjqikwUAGXuuHfXmF3IGlibO+hu7uOlL8yU0EqOyfVul+
c5NHuRRLSOApiLRI+eXhG0o/ZtDYKZPV20NOkBb8EpdOhR7M62hRLNKz/7ifKFseAze00hHP71JS
ROIv/BBFAfF3yRyudX2k8O38Pulc7IE9pKE9ALe6aQusNkYaJdbKkN/ruryu7C/roWX5bEuvwTur
q+DhdXh6ItCHEQoteWpUm6EgNcTMhPTmafW05yVtJM4ZKTkMdb9AvrjBhrR2dzu+NTZaFb9d8JS8
77dIoQPwKDa8KF0kiOwx9M9cCbTIS9CGTCEyb+0Q7jA06O1dvHxmF1EpB8RoCPPzVpliaWXnpbzI
l0LomSNvk5JJDwJG4bcv6KD3E9YfKqZg+6g+kNLTRxcYR2dwMqe/cp6PVqciN1W/AcXDsLe25Gu4
dLzFSOFDNr7LiP3q1WpxFSHCBqQlAMXyLci83Wo6FPzUDFox/x/XuQ3o2fK2bHxH2NIu/e5tucDJ
pygNKYO/113rk1IRd8fEanquitQahu1GFdO+kCv7Bp4oNG9azTyrDfN3TOI6ITpMUij58pBMNEls
jp5iWL9LCxThVIoeNEGxTgd4G3msBCXJN9zQsP2pj6rAawrLdRxa0IJYPZeZopa9Y+X+EaYVHQ7s
I0XbzviUKit4RCwpY3rfL/n2T/UDDtH8BDaDFROZaY39BdxdyeooLpHs8nw79QL6+uhGVOf9bIer
Kauu++gg8DEh/mShB/5NYW4NmpEDGu2f0gEIIcLYDoUINO7Dy29Ts0GDkLwpAFkCTC2kuvlEPsdF
xMoA4fbHbkUFoKuEMn0HBir5cRoqZ3ibP69zMw6xQrmfTiYJSnY8kZN/fets0vTJWSC2aOxZwSOb
ngyHX3ws5+MKiur5Qdhxy0Ct/B7KhuYusUGakwylh8wINwXR60sMigLx/J+taazbDZp0UoAmApn+
UTNMk9ZsCwsyUQBrVZxR3m9ADd66DaB5wgXOWmKewLm36Ggpi3QTPQaBYc4YWHHyuPcIouaDH8Lb
yzBgbgYkKPRIoacTZJsUM1wyNuiOdj1sxlWWsXrQC2axj4eoFkX5luV9K43V4Dcmp9decQXZf7Fq
GGi2pKbQfKATnBIb1mdSekz26n3FSR2nt1XX0u+BpKFwQ0wKjRSe/w2jPk3NsWLgM3OpihQcwRRY
KYlONN6zPn+uC/NEGjDV19C/vqscqg0vwm+DHBaHbExBL+XFgwU9lBQtLRk20GJVRcKqWultwYYK
u3F/w2B4IaOYXrTzXTThFhRYns90zneWvrY7zLjrNJxfOEhRJaBQ1uoKvA9hqNQPS8f9bWUfunOJ
8ChJ25YMEKx4YXkqA3A1x4lDNnslCGVrT+uZOk+of1I+cJdDx/QbynNHNRrsgID29+X1KB6Z4seS
IxQJy1exgIAdtWdVLaTv331rjbkPu6+oHEfU2wi4DETmsQIF6TDPtzzF9tSzZRoT4lWVvhnxXEQy
xjxmILIxdouPRUYgBvmHOOWKT4ofpLKbRAJaOkFrL2TnQ2GY423pLMUbCQDbCmQdDSr+apPNobUO
wNdw70HwPn4aCxFmGvLOPJGFYY1vhAbcoXZ+hbulYia9pgivG4i4XRKMI1axVLskub2OJm2mjHby
kthhJbYqk/zoWmt8TAjHRdCU5HZZ0VV/lbXNW+CXVUSVffa3uWq42aIJkbQkmkW4jVQ3684eVEtQ
onOCYlwgefGH48yO1jbcjYmnhfEFVfoajqeC4yELuZEJRe8vk8kzcZ9p9VobcSwPkqi0vl533/SJ
tunKTJ/RebsXYCqgjCmkBVimaUpTZt7z/icssFF1ThccwTzK5Vw6k/6G84PnQfMsDgUYEOlkGTkV
dnSLE3msvKhqEiQ//hvXWwNlbJh9VobIUKe3zEkcV9h8apq/R3+eIxV3gocCEtOAQH74LGGRTGJW
eoGMQHmEwW1Hwc19SX058blo7jdWjWJNvY4nqvuhxe/I/EHaCtZ8mQETtv9PACZxVvsJWVNtYDIp
JxPSIZWuIIbamfCSxeYmsWRgmVJES3wAx+NlgxDmhTU82/hVeA9nFrCl5xNMeJDSmjS+bfJot5Wz
Iiw4sqT/xpymcAxa1GAKhb180HqOyIAr7f/t+DPoyYzGaIhqtnEpFi2l5GiCaBnDQwMrn7a0+vxF
Upp012iOjZA9UkXA0hz4QzNGUN3stvPmovUmTgYQeUjUuLdNVbYmDdEaGXJIeD20mTBRywxCekvE
wHB4oa6TkHjBx6Hcb4f5QGXeafHm8fp04jc1kwFVYscC1ezXHco1AUfoziczPZYaEaqNbFR9fSzD
ugYO6pBPL/1JEzdW4rIzpFqybDKe6344S2tAPf2JUR5DG6/V2OqAwWVOIEeWGjh9LN39ht8SIn3u
/JnhMWK1nrIv6Ao599KjM5SUdB0ZRkCbpKj4LBlVTM9uFh5LGXh/m9XwdQn/ctPi8cfEemIyDXz5
61XeJNdYXAeGhL6P8xO/OindKVH+9INWb3KcW2TX7A0JPJ8DvFfNj2MplyjSUmJiKmRx4cwDj8BQ
4VjkdUcYskCr0TubfZuN1gDYghfPf3a7iIGWR7NE+xOd4upO62us1hDs21jeS4kqcWDDW6o4G64Q
9SHRtapDOXtZaZz8LCuA4M+w4fZc87+PAr6znE+PClQ4+Pvzs/yGUe5kxyYsiW549+FalKWWHMxR
ZDgxZkYM8JlfmoQpt8tFgRV2dgq9PBd/RhYS+zdo4GX+ruc4tE2/M7hT8CxM8/7FRShtqH8rPK+e
UXtsreNmLiqwjNBlz04Vteufs4Y7pWI0P+aeQIOkfyfZmUID0vu+wQG9mDj8SqPPb6a29pCh4I/C
KIBZ6Ck6IogPW5qCI5fVv5GR7zmbLpN0VFHxiXeyzKOb8qbUiqhbNtZ3ei+L6obIr3FfglJnEIrv
lpS6mv+szaVfVcXlP6/YZvhBeGyu6noExE7XVfQ5Evrb8umPlwvTkSkeWDZB53SVi7tN0mt7cQ+g
nDrInwrPTOUdaagUgpaD0x6F6MvTe9CVXP1oyFRUmZzjhM089ZGq3+CrUbDdlm9oSlhRKLZXz9zR
FM9IKoIfjoFEoE1qSpYzaHQ459uinZ+ksUx3g3PZe/XjLD73TtvPyYGgQr4LWA4wEr5xQvVddk1E
Z0ADLUwBoO00bpHY7b9l8gkVQ+DcttwBitrg771mZVpbnMKHxh4XxCIdG4aHrTWY9Fux6VMlyGrj
K5+roP6qGJK6RRsGkrB+d67YdKM2c9goI5W4ANNLS5GhzX81cYMtWexHhb69vwg3wY3E0GBXI2p/
RnRz2PcC6eJQNTTp2URjELbNyoX+zES9pshhqyUbWYTOhgUYgLvqJcgsN/pevpL9352XqviwTobp
+zrAuiSYn3ADakf/zXV4DCgfp+sZ6TJYGBTss+HkyJeIMEz9vlotmgKSIVrtLp9CHYpX3CIjoqP3
P8HhyYspx2yuhuIJ42+xO3xhl4DOq0Ac+CMp/q1BP4HW5VSWrlczOknyO62VpO3+m8RJnFD8wiWe
ZbYV/XOSwj+1StNRQ90R0xu22O5YJM7Laeaxoe9nJA0+WSuUwk4dNU9Fowz9V64P30dMOMcpSPlk
Qg2iBzkkud4+H9YLfx4FaStZeU1LiRgKHVnvZ3iO+Jinx2rangu0zXB2/XdRUWdBwOuHZuHlLgJE
kLOTJCZqjXQFFZDbqV/D2opxkrl/8ohL5ynSN/ZpnQWvB8G+pg0izZrVWeKit+tCJPy2zIdyw4yU
JCjzlKmGvWwonU8NIrXW6hEiR8hakCOhSeTMAS00Q4DIrT6em/BH6WYr8C7PUbUROWesRCbgz8Rj
zOEcQIDcwSUT0qe75+4wAoR7dr1dDBq+nekMpCLAwFuK+wyi/srwDPATtStcbIRdb8h7CZh1QfAf
HHQYG28YXdY2xhj7Po+aA5NbPR6U6snzqGz6FPGcs/6y+geUVsJJtuKJMHSXnS/WXvJtLeUnWRhJ
S+EX5q8D5qUnU1Y87W1z86F1KJPiIEhNSp1uO1Sm6tuKiJszFssL0sZAJf3yMNgQcWc46aj+niaD
0V4oYDTlVLAZ1RlWpzcvL0XFXv0FRHd3KbywnzBN9MRqwXJqyO4WxY022loJebMObAGjrgK14YUG
uFlzyrUeb3xt9qjkJUUtq0RyC2qEha6gi0CCe8LFlIZjjro8B/uPwiYyNoejDbtN/CFpYI6QdUgl
DO5sFXb2BpX2vZHsHeUngTr9UEVcwLQY02uqx4zDlYONhRcmfFCPXrPGmv3I8HzqI4sTRYKi/M5S
u4rmi9E+z64kAKz/gZSVdDvilRCcMyokWkyoEUu0aKwqGOOLgtubPuNb/1nJ1tqnAXvgdLVCNQz1
sHwgKWxTH2uJejOLroBij7hVilutz3eah9c7z5PqLBB3UHNCpEgqqq6zD74y9sbW/o6Qr6UO8SZv
vUb7I6ECgdwse7WD+6Anq5nDMRwPMauZeKUj0mGGz0lDvoBEhk+htE0rwl0oNy9uodLSkh2bSc9w
Y4nh0P7P7JqSs+yllLTp+3j9ok4Q39at/1DXg/lsyup2aVdIH5HfCozhbklp8VEubAxmevrCA4rP
h/JvSEqaj4Tu36KIBK72/rWp6ME7sP+RXwPSuRghIDbEkXsFbs4KoQd/uZN7qxakhjQNJ08DGOSC
yNaNQTanPfB6MxmrBN4dK10ye3wT2MkFjhJBBjlrGsW3wkuDGZ09qPZYB3kYapa+nxYCnVyJ4H5S
YZWkviZ/guZ+UJX54zfjX3lm6rYtPjTMAX2yjn90fVynmNhP1bODOhLMn2wAhlBisvxQZLF6MjwP
U4YLqyjUTyQWkq4F7JTYmzrMSr3u61f0O8Qwlvw2yCCP11D91x/tXLMghKnUTgWNYNDOWvuFLxoi
5nHTuRNoH37fhu1617eERYx0hGutf0QzKC3rT0P73+I9H7SZGj6ilZncQm+lsr6rKecQPLFSsefB
ZH0aCDXvD1Li/SLJWA73i8Xrv4UefOkvrHB3ssXJnkjyUiyl28hu52XjJXdePXzYkP+Snrz5tFJJ
QevbdSnlZ2Q10tWvf3/zxh+NwyGqv408sBJiOovJawqfpn1AGJCbhloWVBcg2zzc8DhL8WmMveWq
nujFclIKe18nFTSLD/XDq1WKDrfCwemFAgAWMhytNMA3pxTbISuFYPe7sohjMhHioC0cvpdL0uhS
4+ECpQqCuq25yc6snJTua3CKRt8UxRz136rBXXYfwCoL/hrlNKwyFfdzEfBNwfU6FuXtMBaFOX36
Lx7h05cch+SrhBvFuat3ascZjJcZ1kRS5r/uhsSLbDhCKJkBMmkGkFvNBVgHX3A/tf4lhMQkMr8i
DM/GPjFFZE7IkhK1JYjyCmYWkG2KDbwqINf/gmoCTVTKn9/OPSSGFEXxIf4DPOevd0PZEYvhQY52
pqZg7FrkeAXgbSgn+Z5VrBfgbFAnvynqKodkpGx/D2PPAOaf5P4leo73D8yfqZGpL9fnlY80yrgf
gWQn0T3iM97nN5gRGuPCSxCckaq+yrQ9jWxAzhYC70qOBF9I3N+UkCvTd1bFupgS3xdThoqXzAhU
NV5vD5A3cT41yVG05pvCBUs/9FFV7HfVvJg+KGTD1fJr5KQY6aL8DQs6M7alN81kslEYeW8Sort0
Ms2FYnlOmksGZDlofxKqpYiEhy1PuNns0Dt8oukQ252BKcHJ/dQKyZcpO/WREkfa+jBGFWds5UNB
fv4+PcWbzWOKiYCYpiU8b4dn5p8gQ4mXRuNcAtE6QtMeRkOYCg/mHoG47X6RZp36LI+qZatxpiKY
zmmIeP24sqhgSf+5+cbwjMjsvIKiLY+vfHNdKBDcx322X/k65nOCnhyIgrP8DlG0qIO35veUVcTk
olPLaiSG1nQAwXds4aecDCupP7sXUByjUhQK3kPB/4vWcdnBh+4zOP3htoQxs/1sE0Xh2Fy9MV1x
+CxzqhVjJJ0jIrv/Grz+cJfyYABfRC2vts6QCtxxRihxnstLEwgJF0Xia3fA5e6PsIu0dGkhQX8L
yjH6Xb/EfMlsxKPEK8od4TvT6Yrdrd6UeV0HqvtXQTW/qGiyAAKeBWvJRp/saHJ3s49TvY4Mg9Yn
dhhEDbNOGz5tyVUbomYK4SmP66zL309Cjreyxzn+uJ+JPd3Bg9VNBSihzsMSslINVzfrpeohNB2J
cXTdj1kGXrq9Z5zJIzCmLsEXNkBnLKno5t6ZpbVEbpsS/itsjk2CkHg82jv2KRc66HQOuNPRmQHA
Zdb6jwnFG40GGlMgCk0przG9k1ZsVInVr/62SOr2uaSopLBkgZSNBnsjsGfuhBnn19tTeTPAMgG+
CDzRFjrR0PADr8FKWZ9m0Z2RvrUHgmA4j2kgHQZLz/eV1Kuas4cKnb38JQvEG43eEumMBfWhR/vh
IeaWywYhQhkaebXAV6e3u5PLWWwEgc04FtMprWYBpOZ+mKSpKPl4MrFvCa0SKfMHci1cjzfXWVc9
bZUnLXNb4b7z32o04B8pWjnThHfRjaSXnWbaS0wZyE6ReKrIoYa9FFla5QhRo5zXmqIgu0kg5INV
6XU3nD4tEh0NfXdRhNmUDyKln+kSpFhI05SC01VusgMYOkDjtGYLSxoZ6dkczKJNoM8/JLRmbyMZ
1j6dkmHP9YYjquDunlxo2E5v+HKF23XtghKh+3rMHFAv0FXMNl2tcgDegQkBi0NTOtq1qAuJiyYd
ZPtvRdHanryXsO1ZvufBSVyxSqNdgdDh5bZb2Gs+Q0RwhP0Q3TfJFv93uMvvIlJ348QekilbmLht
JG5Kvvj3dnhTyyQm/KMjagZ8xUiUL8P3TVT7pygApHlbXp/GJ43s13kLAmm5XEIHeKi1T0nF8g0v
HPEBHKrwx8YDSGbg6g6vCkdNm2C2ziM245AABJ28nNBr+giOr/XLM4KOErI/jKsa7PtSM0LBceuc
YOy4N8muUsSk1Sfu2SsEZzLO8kmR9ztlY8vyevVoEmsfRIW2U+YrU0bKPIZJz12eABo2AdLRErsj
f4dOGxqMfg0b8oQ+ITvA7k0W6m9qlt/giwRy1BsU5FKFi/f/GkwkLl85zE93PDwY8rGFTPAPvrRh
Zuq4IvBfn9I82/3/Ohma6dsJmZusn0DSqz2xx/lBaqf6VnSxpHu7FxjaZl+4CPMKejrKqt/TbesR
fP9ZtHr9rB8URDGSOjHHKbIy3rjZ2UxSIgR1DzC58JSI3jnxWPqvoLuVR1wHkcjxtzxrxerMinZ8
DkRBFD+5JXZ3nyTXUF0J4rZgqxdyaJPU5wx7L8ruWJMiWscGaqXjXHIlgMBWagN9mZR3YJ7TuWeM
fipGAoZHhXqMwaBxFa3nQKwt6MWo7fq/xw8he7+Iz5ueH4NInOlfdufyMCaX4ZZ+iQNH7HKG1IFo
aRDFrMdst6fewjbD9muvE+U5/pYAcZmeSsLSm3TCO/eBjma28SpKZJp3qR3dHthwqbKa2q/kIwM2
LEZvtG4uRGfXaKABfSCkJGDqeR/6RIP/dUw6YUTuVcQw/XD2EhoPvVCdRf/yAimJUrlvD7NciLmo
BeR6a2j2UVwT9rqSv8b95BxwTxDP+wrLji1V2hwT7ZLgCfvoooFMrR1LxuHV2bDVXD9651tjecZX
cT41DL+tfYNFUsr7thfPoZo606v41WMK49uz3gKX9PwewkHyihN5Rv19jM+0XiUxfGwhjZXRp+HE
3sfIoRfxHG+rnbY4UoJGe2oRGrB/H9dBu3+BsZiUazn0qZLYXKRjnDmA5hJounad533hMgYo5Lq1
7tuQbiffmDFSj68Rf+KwaL4+TjEwaqgGMJBTgwfsucsO7ctWplXHekXNl8yXR5WW+pcyvMsKZQ4m
0PlkDANLb0F+OEbDrtE85wI9MnBJiSajOarXuKMDhCyBZO16NKCSME04AYKExm4u+Z+EFvlZ2i7s
BKYxmgaWUX1Q+9/cuNO8Q+pdZlz10EsKsp1SgkTWNXoeqWtuhGhIMF1Xx8ZyTibUeorAUqPj4cvU
zMemJDQkY1UNAyFa7MXuJ7PFpjAYTQlcJhR5iLKK/DBoLPlYJjpp5r3E5cSUz/+ytV4CP9/N4o3I
oBV7nxWg/PdCUc7gAIkzblA/7dPZPT09jc/A3UkLKJMs0yex4SJsbYGsjsIGf3hEqwAMRN/7irV2
rQxejnfd8VBEhdh9zH+7lXZJQlHcmtV4BRpzylSJcxQyd9pQ1hTtL3RtW5Yp2RWKzW2145yidYmv
WiSyVPZqdz7d+/QFFVenb4HpZ0tAbumDyfCA7Jv0sz8o0F/tpqmunGCwC8RDDMH44iSS+wXufaxt
3pdyF7ktWDQTvADW8wKbpwJhBsxaOmC7pKq0/AdLuKcP6LQxBq+jdqaGUX0tTCdNMMjPICslLYht
NwZVsmPPr6o6AuaB8vvJFVzrMLzcrs7B3MRNjFM4/Ig7GGbV6yz0rEmhz9G5Yim8y1s2Qzt9uSn4
nYvR0ievW9NCV2TAfRks5RsVEx15baXpOFcfJx1suz+gcckVLvkuEaxyC9XGcjk/dlpmD/yxhZt+
8PdxClZg9/WKqB+CIZ+i916WU5WIfKwfZC0WyPjltjMsCNi72m1vvzuUtsPoJPB9oHCUyZXMAR3m
pv1P7LaGNrsN8AOwRcNRcIda61dDvzfq8w97FeXXUTurggNgg3Gyi4mFgjlx0kHzxswsrkEi5adU
FsiYnPJPFqRezYwx/FnJP/3xMA3AY8B+6dOnA8mzgzoW/RPZ2XB18X3LQdkzgbWQmdU4M1UgEynJ
qscbsVxZ90tFi3L8abzyJV2zvTaK3iTwScRYpC3A4CjJiDVpnX6R8V2hhleBIKJdIpwFhnSchUbx
Gza0yQLyq+LJ/d9irkWjIPgU6k8oi/GaWg6XrczLN956jqVoAGiUQ7yWd9u15kbhS4IoGHM941v2
geF8Qe5k8Y81dsW8bC7jDBo3b/qaXepjQ1Fl23TXN3XuFu5J50mCyCgx0vpgxbmtOWVEoDsn2itY
EkZToNTjAV1TTNlP03861qaLYaSuuzk5q3st2dxLjfKZ7c1CN9n6hVC0KRVX5HyGDubhkR41ZtEG
o02xfTbCqxfj04jFH/YkqTNgBmuUqy4S6T4FapXjai8ij3gC5ZxaqgDiR2mLsjsVvoFg0T9STphl
VitUKNeh51wwy9DyzICJO8Ll8otOxMx5t9/5hLDgs1jEXiKr6XEGiuD8rkbnQOWmgkUm6pUxudz1
b/YqTncUP+hDZIGI16+XGYyx+o3RscNTcwoDzTCuOv5RrMe7pe7+JVwtbNyHKcCCtpP6FwroQQ8J
eS5LASoVJPLUWe2DzQrpi4RWNMELmfaqiS0jSl0TbZP58GbQ/v1Nh1MFTwNlidydWrHXzSgPPKoW
jUxIS3ZBT4rhkGI5PRMPMFhXMZCqbjEGUVjY1tFsDRjx4smEz7SW207o0InLZqzCeB3JaK0Wenr3
5n+OMuQEbECRXFx05tfvybUWVXoQEPSyW/Mazsmn7jvXHt5vvry4mkAgd67Jgob3FXD8HR48IBdN
rrDuXFA/dqJaCm5vqDLzrU2eVC7wQZnHNdEdsVZMDgMEz0Pb9MoN2aAq2sDTpkASu4fauLXtuXkt
cbwfnYuVNcahPWmBtMoCg2gDqaLZJRvs+JhTUcQO9F8CIZEn5ggPLmH+Xvl7cUwTPfg2WVtAmzzM
UwETyJAQHTLxys7NmVnq3umZlFliNldIaf/AQ74x+o7ZLax3JnNTy7LPk2UM2zPZTJ/76PukdAig
41z6YEDDUS7618nTrntUWDOjkwB41495Gxa1qaXzBxUSu+vNtLV3IyT+8cmUBxfY9errQAIQGfPX
Nz9IVhixbW4/usAELVq+5mHq47fyyAVf5YBhk89dc2mc1uUHwlNuObsb95FmDc0xqqLcr8m9Slqe
Xy0Fy0Zo5rgn/RAO22CeTWJi33+WFPUW8SctxuxexXw9UZDsPJLU23y4qLTfqgUTyjEzmvAKR4Gd
lKLuLsFHLZhgv0RWGxhkezm1tvOa7GPBr63ecknM8jIYFvsvRlVbaWpLZj2cfS6Q1sNWBx6W8yXk
ryn/nL6CxXvCQzIQ0YRpuuuzGqEnYFovDHBtb/giiqsAii0LAzLLJ6hilkBAhhN8gB7OMWfOeX6o
uVosmh148AjiMPZwZxYTrMclQxj9za2JMEoOPDFwoFBpU+2QUUpq0662ad3nvK/xuCuxHd0eRYfR
uPVPN2UxCD1L7Epk8NBoExGp+QEBjcxZF1JkK5pwBmddcVhqgr4pi/OFNL4iGYRrsR8gXmRT/ptL
WPUQ0MVIuuqjSaShZPktgk7pg6LVyqlr9mKRaFVM6xApm4Ro9R9DcJGjhA0ozEX2yS8FCVVroUsJ
e83GajlMCOa/hvJlNhqa5rkF+j3Y3FDlsg1FyEPO0EW7MxeYJD68hGyFWhLHV8pdGRMsqOs1Gt43
yYIiDD5R+wYnXGFEMLBrvGSsU0V4S0TL9ZBeqhn/FfNJLcMdqzvnH8oCPHPQlElPV6UllSRANZxS
daZRni8w406YQd6TVpjpYM5jMDQLwLTLYyOifZN161kRYqwZrV2cWx5thRAlAJVC6EMtTszkh/Wq
6DtY+vzyGLZNOcyxC2BryFaeC9nnGU+uOS9gEznW4DIK9IL5hLEjrzWnfBJnKodk+GI0U6RpRWIH
0IwSdL5BCEy/zRjU0I3UPC7zedOdO1NtsXtsJFxoxC4CXn8Xi0GdfIMCZEZklqSQNAcvQdog5ZMh
Dy3wQJwM3NL2wLTXZyDC8VH+BbGMaLihJKzX69igTi/viUVBP36Hxyx5VPzRqaq1Ah4X+ZNMaeT8
RizuILHlcS3220WSowO2/FiO/BM2t7SXXT5xdtPZuID7QIrOoBdCXZwTQrvlL2sEmB8PhFDBeZ4Z
n9qhjOaTij4tH6Ws3YOuXyVg2ofcod/QemSafSwQ7eX8KSxiacqDe0+PuBQV8Rn/vJqCevsf4xeO
bzTwTH7B/OF5UZAGs8iIeM9cgDLkMH0ezUB1M6JcCaWhaPeWusT1vfvA0yvHCCqb+ezxTPheoefi
AYC4d0+7qWse/u/eGzbczHIgDlcpmuD6Z3THrRHHkOmB4L4zLO1c6nW55Z1KeGZPX00v5vDLqd2H
HBnnma0r21ugw2jRE2eN/x8oW3fIBDUvpstkmPwjGpCX0UrtqXLVdA7q+GeCisV8pDO4Ov/Ss0Wc
gInZxmzeI/o7wkrqhxzHJ48BEuNt9h0XCNGe56ASKUHWH8vJAgIc7O9c0HgzdlsFV2+kxrKBMZwh
B22KsX2Se1SvEv0J0C/Zl2+ZF4qyzpIFZXz0tfq8U5t5XLbzJXMLnwNXE2oF8Orx61m+KorgTiS7
u8+1yQkMW26VFZbxWCtmWKHn6n+qWVgO+vT6iMku9qgJaxlmMOMO96pcupXHHIDTGNAKmuaVg/wP
vzNOUj9+qJ/N1tZVNP7K5sm78ltfyfxmy0/fEalxg83j9I8wgRY7I8x9ekwlYLgLYRTuUP4epGAD
fG93X+Afh1Bq5vxw2+5MS4ysFOn8x8v57z0tMHN7ADu9LDwGN5MWYpwrndfkpD6VathVYYak5eg6
/mH20g0uDwcSku/ZYgmTVgSQO8lIPxWlVEPEpmPFTJjf8xB1QejXhI9aX+WVwQoaDm3b3khbFZW+
9uFcwOIPdQMTA0/te8nsdkmYKNqPrbNWXOzgbe9eYPw0XOIAXtQd6TOEyGXkirWhduCSMAoVMUqn
WjI8o0EwRIH0ursbizLO5+mPxs/XL1Sj7eiwrnsRUJQ18k5VqjCss3AsGlrzKOQMokURUb47Gw+s
V9Wg+C6yvI8OF3wI5bL9LVbWSKgirnolq6pYiy2P1cJ9Hjd+SIzID/iFPaG6uf4pg7hz2wTbb2oN
+ZTXMX2uOqJEf8h2XKS8Q+S6Em3HIyj9F9XHB0hnRFqj6QYH1gk6Lymj/kXWvRexVEXXgea9Crdm
vtVNaRtmH2FytYVtyl+V3imELPPTqZIEESoo9KzltFugz+f7DFxGdpn2Q9863btIPCXQZokc7V0U
EmPHOY9DGfkS6/3iEi/zUmF78uwgwfxYhSXnVRuIqBSWRsMp9l2iai8egNEPeZreW1Sc8wPmfvqw
9+UTCV9eCquVw9kw7dsgWdT+UG11TnEpUXMlnZivi5/oUTq+0hQAJWOtNnZrCRO3FmXGgda5WBC9
O4uF9/VY0DrloKr5FgljvRXIo92wDQWMm9+HcYd0CAL/5YPFBBBM1/tOBpQ0k0gQeCZbmOqCnuCH
l2QTXHqjYlb/0yQs7P9eYtTWPpSKN5kk9Ebbxla+vaOe7WKTEOJWHD1fZsI7yURqpWHBSiiuKK1F
MoMvEhNbSZdoApzJCzEaLj0CGcGNESdm33hnaIF7hFn57SNDIRBa3yxpYHlJY/Kl6DaHMmVg7Dre
88WFhXqX1mWWfbSHSwYNner3iCr4SdHeFU6Wk0EH/mp/98EtGsqEloNMp8AsMEoN33SIirImQQQN
SbfvESU3DX/K0ZrxH+PBJMbaHw7YJyTnquilm9r3maoBFUQV3vNG9cQ1cwm+LenjA/02ksX0X7Im
qTT6ORIJwP64cvQWLLwHH1C3c6Wtcrr4Pu2eMhf2Ux5J3cHXcImrjSalCTIdYONJJWDm3SP4x8AX
zJcER5pUQgHtOl7jgQt3Q0CBAtfcrP25fgiVZckQnJrRUzmqFMT60SojPT1nOAvm7Uh1B37qnpAz
gZu77sbcc59xIBX1MtbTs1SwuNgKg8C82xBBlWxpKIoeuk97v8fU8WjiLVXAENfgmHQlrXAP1HGE
ke6FXXfsW1wRzolxGBJFQTjcsHCUTqU2AghvI928Jq6dI0iuOa1wHpVHjmhJLoRWYLDKGKCC8OTG
cnSqHpJQxGGnGouwTX9Pa9EVGR2XMWokG0D0xFyChvQY4e5u7j/ZS7i+nQ9vu+6vaGUyfZ8Jd/lm
LqJTOihXBiDLJ283TYLO4Ui4YfIYMfVa0iN4zDR/NlKX0z3Qi74F61au70ZzoXhwIMKS0L9nu+NR
rNgPm8ozP5XbveF+K46KjRfepWz+rTV8qC3nH5j644lHmpWI88g0go7nB9UK1seNbZHrRsgB8dc7
v5UKilIVWyCJxDVpAnSH6cgkHxN/SZsU6wi7OUIRGPsT3nVx1ifpdLadw9E6xs0RKfUkprNgsZdw
70pK3sO3dMKvrXBGi9lQ9xSMygSeZVKiZNAqAm4LXPYbTj53pag3e3/PPpyIfCoMpoS5ryAWY/bI
64Vdewr+Gv8JxFNsacdAyhfZYcakDQCltPkiXiIgTox5IokydSqAiaktvIPuDVxPj6TatY+q4A8M
2LwUHeZ/88pmba9DsnPTXSHtdE/VwUrqLmWq+UHd4hNI8hERqJfmNsRSJawm2r1fK4Rs7NrjMg+S
yoBOTZNKLU2+Ts+KHmvWh5fMSnRf+wMGAxFrQE//IhZbno0vEjYlREJ0HI2pi7rjEg7Gl4BcfXDy
hgclERNEh+kkhrWRSeeJfdA8tXnGli48SJ6eOPYfe99sfkcfe1PPLh5IoYrk7Mcc658McmjW4gip
Is2s4m4gWSmvRywZ6tL3G6jOZ2lT2FIq/e2N/iNqxvA3EOMPQEH3rzV+6HAgahNvA6yi6mxRyQgW
gS6UIPZ/6ZKQTgp27JESbbpRc361qsL/W1Q9fZGxPQjDNMzcX2rg6E+eehJbwuPfiLKRSbh2qb1l
pajXHkTuYMjdqGxiltQVFqsrWXFBUgFarIVH+b6lmIi31wbakCaSeen00x+qdFpN6U9ZphP4V5OJ
ecltwe5iwgkQyUsTFzDvbc/1GSWulwqXqYWNDfKXu30QwVV0m+KixsekoQ2PBiujwogKNapjpGFd
L/B79aLBK2y5w4y3IXOmJK28/arTjJCTy4ZPL4+VPvOL2pHLTn8gL+5X5y/RlKkEVriIqn0FqnR+
9RLfA31dWpXAfnGWfymvJ6rjP5xk68REkzYbOQSdbT2llzVk3ZZb+FY+Iq+EiMWUL45631tM9i+w
NyaV7sokpVbAkIRUKRqVG4ltKQT9Elg+allHO3eHLb6355cFmuKxxMeCvz9W/ZRhJrlO+O+3Oclf
H/HNObDEJ+Kmsv8KMDo9m4vjdzOhOnmFx3ffzqdph1txSfT0vhk+n3MpGIcQLijMa6UirRKLMT82
KADikQv4Z7/IBRF3It84gkWBWRuwFovDWqB4F9UguABWvtU4lb2XzkvJ/YYsJ2n43qPT6VSDjMW/
uOzqbvhjfmO3C3s/byHYllWtl2Yr/rgOlXr/ieG+rqi0q5Dr9iUQIfjkPAKlxdLY+V2oBkXO6FA6
wQYpGgryRaUY5NlN7ewbfaoYNc/TohBzblgAlppT9492Akj0XGPUJWt0P6vGr/5RvyGy1qVT6QPU
mRf72OAB84+3Bg/iDTJxuMYYgM3fnkHKaB3mD8JPFklSeLo5TD3KXTdDwoqVmG1ns5lU+QvSPkwd
UNEdIVmd8lcJFHmE+sMDOfoq9Rsr668Oj0Gp5k5Auv9Rc7zQQWmPcirQzU1Cl2wlDQ+KU01lZ4A3
QkGQEkh8CoyBQepuIXwTI5+7VC3A7nbDcy4eQ2bkW/+TAS4DeLvGUCiQAbQbwqsEqwYFiKoD6Baq
1NiJmfW9oT6JK/rCY3SocZ5TRq4vJhlQPHkFca6y+CQtJM00ofQ3GKqrSP6QXCsbBcBERpNrpTC9
Ly5lWIp+bv/DJMz3TB7sumXwE4++jNx489QTeUQOItzZN2pQdbS6WxurjZbyPzIQcbgJ/BacRp+2
MKdIwKpEVN/Bg2Xi4ocWRlhfZq5Xl23J6Ld6s2iSXx+y5zfnkDT67+caMLlUn+vbd05mRxRf5WnU
K7X96dZSL0OwVdFFFlfF43wER65MDD2jC2ZvVrKMOB7om96r9mL/h2HtK9hjiVm1poCkcQ83mYid
x1burLu2l1SXglfZDPx/slAbES6S7cR/buMzsDYltCORcAIEYLkc+V4xB0fx0t4ygBLXzzX3WMTW
E3G2F+vvKQOPawIwVRrwxbBHy8U7JzmSjBsaBBHbrP0MY6Oie1mTuSsMfUzh9d73WXp94dOIAP7u
zdlN77uAf3rot5hzjppX7wKJW9pVm2O1A6vD0xc3PUykSoNVSlHCOoKCXicD5UfvkB/H6SHP7J72
OQPszOiCFGNLmSIUWdZ8SBMmLde1Vvt0/tB4eG6Mriu3BXjZjDpyihv8rp2TsC4QXmLS4Mqok4gu
9l5EGsVmwlvSbhvUJFtPNnfYWcrLahAYzbSbOnh1jJHy4oOsJIF4Y6KZj3FUnTHNnNVdAQ03DstN
fo2MQYopjgUKNg629vy51Z3Zr025xo2voCJYt0GxtEX6AnUar+7iDForWUa42eukeH3VqAfz4xp+
+iYCAKFyt3GkoGlE3UStb53LCZlUUTrzMOITpNKtzFMk6R+E68vhUTIPb20EzRSc3MaNEzf3DmyS
mAkBK/52TLfXvvtfQTNSjfNPtrK9ppPWJ5By3ACHKV/R3+JlNO6dYBDDNXn8dBGJ1tKQum8tgYyK
vk3hSQ2F3leB0tRFFu1Xjpj2Hsc+sOeBotKaTWkzA9ghVnORacLTeJhsj5dOjn+7XJFeYh5cGiF/
NWRnyI8UMMqPc48SuT79DwwIzmrFT1wFzZxXFn/Sq7Wd3dpPD6U+iAmLpvYE3gBxz7iPh5Y2JnJt
RzCS27sHgxhAtwT/iIa7Ftas09I8b3sHWR6kiVchrQ7kzJuyAWUYv+wlYGdjydRUP+mb4YWyEKgw
SSruJDZCAT/f9QNJuDD8bMzlGjL1oqvpE0w6XM27R0uiIl0Zctj4kCQKa0xboEOLNNSZrZ9a3Ha1
ACIsRQP3Idut9UYemxtxp8SK9bokXEsLUzYYLB401amr7ldUxO7bB8qZEuyI5vaqRBluEQY/N1zZ
8nJDjLx4Su52oA0vuCpiDm7J/kfP9HarxerYOF6agkxYCweqbRpyuAU8Udq6H9cZ3BWhDDg0Yyjg
YI/7/6pZ6tOQj7agcG93mzoFzk6aey8hJyRi/TlTNs4jGdWsekv/t6WykEMI0nn4DggNjyPoPXRo
uCWr0qZtHZxheyTil+Vsf+ZD27tWO2wT4h4qB4gk5G7e6olY9BNmQVO7ZzQW4tHxcFuTaSA85w3V
+V/QeG7Ii4WI6LahYrNuFxmApNpnS4jxqqAgAADIxNp39bGnGvpsuCCff9LX7UrP2KT44apkTV+Z
rx/P1yWJ0zwl9N0gGiauXx32bJTNOar+CAOju787yFXOGQ3mOndyb0l9EyGk4iwblhxWzhwupOvp
bwNIYtJ0B5OFhpE+p97Kh3BMajZY7T8ze5nx3deCtIwyL0pAxHyd7cFGLDv6f3eDDM+cKjhAywWs
WPrNMqayWTN/2/UUCbtR9lu8fg5Y0jLPN3YDDMVdyYkES0wU6zBWNWR2tJBHs+zZ7Dcq3STaHF90
6hzTyHdncUxOSO6b63q1DIWL8yVMnlN0TAHVoLQHZ9TPoBgQ1ibeM4xS9gTJg59QJzsfEphK5Yx/
1s+67Ms/EzxMZTrWmKRGKghi5Xf07+YyZV3B6zzEJ+dFTlkSKLumAFc5qsLk2KgNNxcuQbxta2UT
TeuR8zLASIg/zCJ/JrvOIuN5gesLv6QO6eE8te3iwyWDAnAyfIQ0FNC8lxikr9p3uCcPng/ZyKNy
RSnMqQL/In2z8QyRx5OueR0Z3n5j/RtslEbM3O0RV0A4ntP6OmI3ZHM6p0NhP9TsOL2YnBNm0n7W
hdk9eZDJH64XnYPRcyhbWUilxTfLsSKa2S+9/dCt8AUFjeWVBhFtZ0pOyLTKa9k+HmLl4elnuZll
dLVMrbhX9Et87yQ3SDgVi0PAs7MCdXFBu8Y5xKl7KT4iPrNi8I7sjOEMLSmWtuWs/3gAkaRIBy+d
WwNpxw3666HjLuSs+gcJOpoCa76fWxwdR8DuUK4xdsF6xQVibuqV4zD8UlwmXWMKf+zFVC4NG4Qe
eF3Y08J6s3SThu0PMR8CDjEBqB3QPfhrXoWeQjjCClX0XJ5zjpV0f+3E6AsGg3cqPuPt9VsIshD4
yAwCrD8rUDbzDNUA3/hlUT1hLRx1eWErnOfcnB823dFve9WFjwfqyjWy1zA/13Bplh+om9sOMKm/
xCXonMDiZ4n8cVT245BGD2M8jfCNPiA8GG8NGQqH+mmQe6ZZp9VpqzKURPqWzSYuVuSawCTyjGuX
SbMO/TCRGH7KVHrxiJhJbFzh++nkB8luynIDKYB7Gn+IOtIQFZQ+o8LWtDQ+SIPRZj8RQx2cMP86
ODaJ3S9Uc/PnROfoAx/PtaNTdwRih9nfFVGX7JBK93FIO428GqnYzXUE8SmGpofTP4VM4qC62oSe
nzE75/idwKZfb9hRH5A3PrF/P3qs+ydB7zp5xRrzb/CERab2hQcc+vTKYGACZa/6xWEK065o5gwE
9RBmqVR0Cm0iYjW81WU6mX1kbzlNaRocf28kuE9j8ilEfHR1XuX8VODEojlfVPQ0aqQ8dfuXq5EO
ZJcEnYI2ShAIlO9pfweeLGBV4S/MXRcIrXe4PS4E7iRA/syf+A8CJTWlHDxmufmtRj1UpCISnyOA
IhtMPffjAnJ754lniLZSLotYGmk163VHS+VQkIEwH3VAE1UHDSB5Ac3+vTpEFrtRCKtRKaLQOWXE
t8F4IaeVvVoEzZhyZH3x3sfMoY+ZxKQgBPAPn9rU+Fq03X4FOBp31xa3tiqQD5NYOYr5QVsRw+jT
VX5zGcrHppr47H15TucRL4wUIk8jhw8uTVoAkT693PJGwRTXhw+gJWEkzwqkIFqV8yakZfFBTbFW
SefK8QDrd0dEhZ6qbqtuaff3VB3ym5s4SXvLPo4MPp4ApjERCXCtr37vbOjeptfkPAEVYXnicdzi
wIMnnEtXq9x2fj/JqOhoFVseltMyBvcHIWngSO9zwFzaxgn5d6x/cm5AQMcLvB4cOoc1dHEMnn4P
Hcvz7KNu62axoamWA0ubhP/0CbwKKvU+HYtKJsMbwXZ8KJaAFqaxOI8j7ZNbbZ5SD2KQNtsGg3w/
oJBMPzGLvY8g2V1umzuq42nyjPqDRkKuCdJntrdOI2SfsdTui5CtNaNL+eicr/NqQXzpHRdvm9ts
OMbq9rfk6y/ajy8HwDV+hG0h+Er+O6efaetPjBZg8T5rPD9g2aZssy7ZwziiBo0l8s2WwRK9Eb1I
jEqYFbELe/OI5Mv+0zNeTtemBO0A0mIDkdHZ21v7fSUNgn3H7mCUtrkcmTqaXMkYdwC+Z6mn6GOG
giF9Z9fQ1gnOA+FdhvEts2qtAdB11YpKv1lQgh+7LK2QKEYbSsEaGI/f2Qzq56p9pz9czo1iN+Cd
ONLd1t/is/0FMoJutzTImaRq6y7Z+hB4EO6CSeFksJZwoSC766M36l3PO7fi7QnXzl7mn+x1Hu4s
ljhcjFaIvM/XbamShn0Wa/qwQxx3IAEW6jewFRcA7p78HPERr0X3Ob6ebeHNszLBFWwdl5sq/Fsc
ACN8Qqcusd/aeJU9qTcUcaIl783Z/1iF3UMM8Gih7bjstCHTtX5V4h7aWm3yO46659sxkcZ01r48
YyooNZEslAyH70hPBa1QMi7p1eWsDKuXu3tVi1ozSKEAzzpVimzLFRep8uXeYMT6x9wTaPiDErnS
M8CBVzCncvq+hUL8cLGT6cN3J3X8RD2HnpqyyB3lQhb03pdrQMCqVuydQfTWjdH5YXrgy60ITZyn
xXqWUNGDizWelG+ngfmMkJ619z2RE0VOnsZqqb3mQ97vgYA5cQuaW0Xb8rvnzgUBunF1ta8smZOk
/1UfZ9DFqJrHagjeXam6VxT0jcGoqCHm17DfRzRDxjJ4b0TKuTS+R5oftNWscJen0Q7N3R4J3OHO
Ys1UGaWY0EZOxXSCprz4oXtxObjE6ih94mNLONUuLtdZ+5bQF/uoGwtGwJ14LUgedyp6hfg1Kf4Y
4R8jRiihPfAcEyF2VQ/ISiHxW4pDv5o/Tw+L7yBBc7OMSsZZBCbFChVV4ol20vmS1n5T2l4f3SfZ
/j2k9Mk8nd7KiHQ0EP4K8n0K3FnFTs6m0qvt/4WjsdgIYgDr4JuzB4yhRMTH0bgWtrB9olqZyGmM
UBllnj7DctwZaBWQvskwZXijgc1xlE9vSCOxwEwSIUhxf6NeJIwCNPrAErS7UC0YYyZ3KYvGCOHM
YEp/cFdoNmyJ3I4iQNmDZ6mwN3x12d1o5iM8InWhr9DwOh2UXjdrA+9VKp+B3zsRTFWduxhItma2
Coz77TjQIjn1/YT8ZZ2OVTNzG6MUZjHxAcNAFyYT1hfLEfZD6oZGi/DPC2ntsHYyZ5q7bPilTxRQ
YxOwSyGl9HEm4WQVBMMdS8BIKSWur1ub/XbpQgx5FDORFWlBQWZOaMwdzGnerppc3PY7VvHlecKL
kdg3vURVR7mPGyxLXcP4eY9YNQJUXJFO38GvehLjKi+rqq2NrnVcxySQ7EyYXuRhCsaIdZ+2oXDz
gavGKHMnbNurC68b8KFww5jIDCLC2KapViRW22nlOy827RM8itnhMPKFQTNmjn5FIYJ2evPQtpJb
GGhd9wI83gk96M+vHPwFS2h9/OP9OsrVDA5wl2yhbKrM4xgK8MWQL/KbWjQvpACMFYks8gy3nEcj
Q1W1HoRsWBsFzcA5iIOsok/mpKCxmd2krEpdd2hKcjPgiaiVEL1bYCypWIoFAFUKEz544Rfv1TpA
CcBtNMApL+Fw6uOyq4UyGkgA12DpBUA+TODUeAbW0w7cBNGctr9koEEmJXGFzcKZtysOticcNWMi
sAW2seb+l6XQhDu8i6ydw4OPD3ZVrnEbd+zVkE7j4EvlC8PH5cgH6EOpVA/6AvOpmMzglu1iUH0W
bxk+wqvEShEG68/IHAnGCdvaSwLI8cRPShOwAm/k6n0s3WBWmDhpMEWOjd+THyNehPw9eINT/UK2
YA+Zxl+grhHMvlWcRHKpjre03qI7RcDUsDg2dikqBzixD/QQUAcxuYM0xE+XiGXMgl1ooZNWhuWQ
UDj9gpTdoft5OyoxVScDjPT6w4WVgxhdYUpKEx571DOjNG4sA+sC2vgR75BPaY7TGqOq94kxSrZZ
4BcN9K+n4j3q8iiRCOSXNnCDhychy3mktfp2VMlNcl4b1Ygy2JbnhkYnrU5jqiwQKk0Kq22Dngc5
pcFkPJ1NsDFmDgq48Uhjh9S+BZ8LCokHv7WrXOapYW8/skpCgO2bg8aSIh/5k4trAt0RSAS858Wa
sP8Sv3ad/gN7Susg2CYHgfmlFhQ9ACE+eQ68MTrCHZzJJIKIDFviI5H1opOBdSRXlV+yCFCivbdr
D3sRe4qYp1evV8PyxAK11EKcjpiXqNAMyy5O1E4ItyvHz/BY9pDqglt13NxZCqFVREGH72udOxYe
lBjQMwBL3pubKeunlBFef9eNefHSNLAKY3it4UEMsK4xCZYzYT1yv1TnJeVpGzomCW6q9CXDjBcE
2kuoixALghJt1N1zZgcBGQ3qEFqWTSVHwyyPPPNJ6a41qg7KrEZpXonSNC0JhjUKuhsAmrcDwsVv
hq/kh/CCVuuLt2uEfOF2vOntkXOjAqOf/9Smk3LpOLBKemaCmrIqP95AKuUHaNw92/iuXBIJs2sC
w9YE4pVkOphPHoxy2pEaDOgVYK++AgN6wPlXgvdyTpRLTgmNdQ01B/qraVdpw0dH7Cvb71Pkdef9
ldoNcjU4W1v9MlfpfEpiEmc7VFREyUSuGCe7rlFp12q94AOYGKxdiqstB/7oisO+sM5LPnPTNgFF
GYZbQemEtFJ9bd5q6jWEdqW6WSsWaLBSNkHDvyE/8DdplNulVCet7wz43tm3kckTVXzREAxAkana
rz3gIFDD/zpfjIK9CICbeaTqUfxyFnWwlhgrzkCh68nC0OmMKaTRDokqjpE5GGL2asswlBi3jVq4
FyiplSUrYu/jUyqJZEfwB25nknazHy2gWp87qDy7p7+oER0aRNu3Px55JBDdEAUPXieRhFeowNk2
zBIr+szdKwYxA+fkpXI3yKZSn+4I+e52HXaV6ubu2iKitboO8syGr0VrTmEDnXSxD2HZgmBSVO0g
+jipPlKuGRSKcKZCe7vRSydBESu3l/Jt5q+iPUIfdTECI82aoLQNYqX8drNxvp/f/Dc0wyF7ykMR
+qsjBTbASIU8FZ6vBtKjX4IAKbaPfDaVxwwJEPkT04eox3lOxVMS7Gd7lsaFpmBVYG6zecpNdQlk
1zudfKVzkVKbgIqAndERPzPTapqOX3xFAr2z6yj30ExunOZWGTWm/b/uWl/RGRumJxcXIgQ3rdcu
qEnnHD8wsAiU1e4KkoKvW1n5a/Jw4N1VlXLN3+Fov+9xCTRTahtSpbTbMKVH8h/2HMA5o9jOGTRb
MuSpBkoXtlf4D6RMfRfvnKnUCv+025j1lMZg3nA38zTrG9K5tAkaEU8psBpLTJhQ4qTcXcbXZOeL
1dsx+VFGPLHqcoJRAEuGsdHiGbxSKUfJE/sA4Bn0H6aMRx9bTRCty5K8o0R2oJA+xCSBLkjmh2G+
wuQqryqkV31g8AZ6bsrT5N3lfwXGpiJfhuBcUzxdSfZMIq60EyW0NtbUeAppgeClKAeZ9YdzhHxG
2XyAma9+8WGgTEJQbzRhPfwm36abqhK28wNw4rBjoZTe/PayW0o153O7aESsYYa1ZUizccAlZt6l
OzyKWo4iRD+H8CIFK0Pj0HEJgFhJS8NrhRsWX8S3JQ7KuQeXCkpFOiuO1EdAlnaCgdaKnJSlpcsR
s9b7A8FYtoKMFhbbg1DAydYMoPa7iaUqAvPAPI7q0XoTq4dzJ8giOLkuciqYFt9zvKIFcwYPmNDU
xaKu1DZ1A2zqllOnaKFMJ4GjkRGquOp0tq2X7TaqTSP2V9y/FOT9tyMT9mr9pgNbOcIoevDnXE6B
F59MrHf2OhCimwKaq9H3lNnsYbp6Y7yRBmiBCdrhTMuU6WM6BVsarSfortlpw20Z53mzkuXFmrdG
0qx3Ofhy3Ri8LmkkjwoUcHDE6QQzh6DragT5Hd4KF0d/BoxxIR1o7tekhZB29rq9pnY0KhCuaB4w
Znd6QsfAECs/SCbkK1M1+9E83mHppGz3vV8lnB9MGRNF2+2cITMiI1VKoosEK/jzDITLobQ5LlWj
ZC1yeQUpws2kdHyEqaoWLIH42GjTLqPTJLmbPvpQsBUv4kOunjNJXjKhOvDIYV+Mwohoe5FBnszu
3xmLy1Jk6r2mBnTExNzyeiUN+LGyz1lo66ZJLY9Rlrq///dWMTwlx34oOAbLaEQGSUGsO/BDGF9l
MYUmdh+qg7Zk5eQrxS2zjgZO2X6bL7kF3+pv7cjes61lpZC7JdQMd9MwjGju9dy7ABjy9DscegW2
u+UhXrKdPXy3o57F/D9y6jAU7KDCqdMIyLryxuuN1dOKVKlhTuf1d6WLpNniTXijAIRpF/X12lza
iq5LtZVbvCjjSYNcb+xY0I4liviAiUY8ohQE1J60GqkOgE4lixU3cdZI7zFkPwMwoLdk7nghLcWE
iqy2+/DN3IBFfZGHPjEHzKO88x7Kl8jDumI0fEc+IIApuvIg6VXdAYddA4IlwQqp27vmC7tWQLwZ
/cZ2YEueyKk5cbcqnpuF7or9QJla1zTLOCnd+gNnEsjVTv9CeC734zSL6yS4grnwTSavoiguJAOK
MXWs8HLpN7ErfIsQu0I+OlmFSR8OvXx4Tgw9NsjvM6FZ4Ii1Qmvt01Lu8K9KIQFR7cvGdNiLabC+
7HtyFbhbwsBi9HXUmHbOBmZeEXv6ByLFioLxsPod45L/oqMbggbiqnju8bvk5Vbf9Ok+x4vbcL5R
t3Hsp2AHO7X92bAZugTMujE25hpSwL/h6363v8rSfLk1rANzsPe9IDQnbQECmbFn1Qk6hY2a1cVA
fbo3rEtUBguaDYeBEXejHsugwNCeuUTZb/g3TcHm1hlKv+NLG1qJqlmc0hTNucOZ5zg7LkFI9oab
QZIEpgCacUye9kWWAbkhZ8Pk5nw4cgynTZsG35fQ2ThohtnAcK+n7liehEs2UU0AiE8Fi+AdEqq8
RweJSpAuDKjY/tRZH9YX9vpFbmyiljUtUe4Uel5Ay0XxIl9AX7Ucg+O8cnz6hJM9ry9MjC6PRJwq
OdufO8umOSxP048z047BuJOhwGHPRKSP70idzcdYfshco0/GtmaEzUtvOCVXpHfUkDNe8BoHw9Vr
SdSbIBneEP0nmDsgxR6nH8Dzti3RX3T61flGmQwIMj/87Ve9LT7+aI2HKRVziyTG3C1jf48fvyAm
9pzCVTeUw6CiW6Hri0E3XMa0KonPrW4CbyMr+rJu1aCq8MwX7CoQafncKIkcDhciS4uY17q94h1S
w0lRV4CvUi6iqZog+HbHmFUkAPm3R16FCOH05LrVGs9fJ/4PrQXmwsqFVfM+fyCNpHwwyctgLcVm
pfNE2vGBhiIcHLbm99Tp7uwBjRk1jufPO5lU2YppvDUljQqJkIX2ZUn16fbuPHwltte7qBlfBrTG
BdyVk9MTZ9NKZS1ZwAk941X3MTu2TLXXr5M1TrUVTj7dvB1/unYod8cq6iQ7NHvyUnj3wuTVvU4f
50jBhBAEnYQtBaW4gLVtvdZ60G/0xk843n9WjTu0APGkEsxAfHy2E9pEQOKfBSsnME5gif3kkCUp
9EM7edqCoMND6W/PqoNQZ9SGajrG2eaUURyeF4wa3RxclrzrwSAtItBPjjEAOG4BxnGAvjlUZz44
FLBOoKXHNTYpNV2WJulvIK72PnUhXgJv69OqpYg+dzRFeBhM6Bmlbnyw53CVmbyXokWcdIz0WeDi
LkXtfW8/Vjgy1UklRdAu6wr8uw+d3aqkbnZUDEPr8/cUuqCncDJQQc+M3DAzdRxREOdVGt0ZxrdN
uqZFc0SnPFpH+Vyng/EycxzYJxLHbLe1no66HqFamXqGdB6b0LLBHBGyGJ+PY0B2U6Ywk6rYCkAF
39JRaQdh+Zmdyokm3wc/cP9UxyVv4gJ9rANL9D5mMgEpOPFsiSvIKuZjWtWW+KsD8L5XrbAqt3c8
IjoJdvNq7eJZKNrZx3+CT4YILsqYKf6tse92pg7/JYj03soDqh1a/gmTDk7HBlg2BeQ/QLXiD5m0
l8TiyeTZs6I84iAENzjYEl/t4T/bnxdM5UBIOlytB3v8VJxQ/yuLoDZbh4ZXdNz5LXMPZImhKVOt
a+bXw4fcM6BXg/26YIgB7wrG7u8kAX9PZ37lv+NHjeTQbhQ2Os+18kNyBBuzXzogfbRhj5ufL4Bd
dlU+S8tOsJLbeIqDcRGDhfPr9O48BX0iPHEivEQhV6s2aGyEe645I7z034ILfSGHExN0aE1tuhQr
9gLXgtCp8+hgOueRZPoRz4bXw0K3BTpHIj89hnAGyl9pH2uk6hQRT3yatsbAIuLHUNXlTDu4SAEN
HxsmBzSN38REDRAgD69RqI97iRKce3tO2fyBk4lFbN/X/rA5wPTFzmMUg8P4qaNQmTwWB4PfOtcr
KxBIxJFS7MBR2NBc2v5m7pGPDnXC4ZorgJfrCAqAAFh1Nl8dUYvrMBwUkdIkMtmtCxdJ8jVG/Ppl
2jj59CtLmB9F/DCKa9y/dlHi2eePhFbHIQWcM5w1Yp9aDdTas8GxHrY5Yljnx/2hGOMZZDcM+ko8
7CmHaiZGNuy3WppmQ2GAotbif46GCE05HCECEL6eXaTpvL2CSmh2cSRC9vCXEp4oOMmiO0nthx0W
nyEy09DHZye/Oor86Tx9QehIHBhV/X83wlqDR40Ys6nPbZvo2BB+FNvTKEMK+ujEecP/DPIEO2oM
rPj+DZWG/nAq9wgVmYqinm7hbIEcWjjc9dmA32ZThfQgmrHJ8hWkVz0gvJHZPuFGbm3rBmY2cfTC
MoGDco0SNDaaA1ZL5PMgLPphLJlJNyzvRggsecbJeYwNAScZCG/VO5FxICZAGFE+MFNCyEHF2HJ4
uj7lH99dNIuLI06bvC1Fu7ZCELF9mHGVKn2Tpn03CBwR0I8iz77eQIGLpdE6w0DnFwyOyujGaC9f
j2mFNLc+g2oOvSy6parnvBXMCLVSCNaccq+/5fcwcygSQw03E+iM7F1oErLIrN8KyFSQqFZOcZmS
JAQp1UKv7fjYbLTnBjbs5PWQRv11XvfJtzOafAHhUNJ1bJ7xuqoQhy7JZF5g84Z6m0/gYd+sC0+E
EjTb4vd8gHFCWyypIxP0vz4rNkD0O7qMVZntYv5qHHeQKQOQW4LvwRnirnexdApsVjHZXPpQ1fJx
4mSDE+QKdLoy/sUkNJWTEQhzZh3iJHS05ZoCwFSDaHUwWqFx+LieKgsN8rA/UWm1aHqAZ+jNVFR+
/Q3Kcj4JwT8dS17hzDD6mAh//ZiNare5+2FlUtzurUnePMMMK8If4S8rcjNzl9dBHGVFm6BzyxPl
rpo459MjCS4A8S+twqtoJUHnL4zWFhkgcZFRSuynGSVfl6k4b5XTWJtP8V7n0h7If2IzRbZ/KQye
wRjJeDZYt3ZyEn9kYBXopiS9dAxZXmGu1LeDUxabsD/lT/BWEHRF3tBXYK8xOGm+EuZrdOTEmQS4
7mCmihA0SA6T6Zv1inw2XqWYS/Hpj3b6DeJ1NjTl84q5X/YiAqhAUHuB93lxAKwt/8KxzL71KPSB
JtufJmx15iPunM5gLrOV8QgMnIgn061W5PHMNPRroRv1l8VxIE+ecdMRPwwL1mI9lWuvOTYRzlCP
aR811tY7TbN7fHybDjYRduMARGgOxd34S+BZQZII3xk7nE2LZmJqpc6IY+XSc8Zt0bC1sNY+rg8J
40JIRqM533OGBv0IoQ3zc9ul1v2tCaPX8VMSre94UjIrnwGNAdydL5ndNaVZPsOMsfZcmwPNvkB/
f4VOsBm8E+ZFrE9hIBDfPrF7yhGb5CqU0Po//bjd82tzhvddW6TXnQRzCbB8U93S4MK2gu5s+ax5
4vSNT5yRHc+4qPJUeSjUZnEL2xtb0m7PS6u58XYL07FnfGoN2fx1ME+0b3ye3qXgJLFh8/FvcijF
jKVCgAbSwofRTAo6ocQ4p0hsZiezTGHe9FImfjCNB8Uw+VHtZk7ZVi/JyKKYzxLp7WSXpalF1Tqv
y/pcEAhQqKmfg+I4y3RiFQYafdnx71yKzuy0kzcoBJ3MpcOffG1kXTkU/UBTWBg4XFMbbTzCKPau
o0+Ojf9uxRBDnqfg7Vd7jo4sbRyqQZIEIP+sd2DNMmIfKRXT4DvQRbYiOHWeaSHhEaPWdB71SoCa
bpR98VrOjFZcko/0kqqjaqZiuAqlP7SGBVbGS92DcWH2fPqjBEwTrKdqM2Qysy5NLySNFeMIbXAD
Eznx7t7JzHBfx+Dh5wxQM49ccPUw9BAxcJnKfrPxwlMp7fBC8q6CrlHZXf5poVN2H88Lhc2eDQe/
4qVq+GuYdNvmdZ+6PZHwAzf10gMm6pvF4MF35vhnW9ejWC06pimUH/KiuLarX0nCodTsydXM4Zy+
qZuaxgVLo+Avv/XjTX+DDzttIubb8Rp5C+nyvskRXbfMB9hW3/pOY+WuFaJNppmJo9oS6AQp3Sw1
kjoVgO7SyTIBwyhkSml5LqU/YpxpNkx4MmpOPKTyoaMow4D/w+tFmMZS4ghLQkdEQur0pxW36KYg
pxZCQSIdWP1omv5ViD5p2fULUNaYIu63Hc3EJ8N736bajaxngoKNuRTrODq70kCeL5v+av60eTH4
WrmVvZzHdGdeViiFnfwJh1Kp+IwtbbpBmqL8/1t4LmRF9LIryuNUdJD892QlaDlrrwSFR/HFviML
DrPZT/MNslw+HGYlWODZr6mw/KmPHbX0GpmkHbIefH2TpVZeSJnGP5Pjv1yxJGXhhWVq2jLpy76P
86g0x39a9/TN+rJM2KiaIeofsjhs8D1YWPfWYqxfO6rR81nyuNhB0ViWC/ojFPHpgtOH6nBIBV6u
fn7NHGAiKLQaaRzaNokCR9qgJL7nfKkjucqYsn+cvygMzPhcPsbcxvXgoNqBoG48AEs+8xyMVEle
ArPymAQarZ9DSJhGzk0ASgZoEYtCu/0+ynZMQayFIO4c+r2oAgFRLs+dD5tHY2kBc98TYGhrD4rd
fNsCUk0gVL4RyGUfNcHgBrA2cbyEzaac0BRqoHuQm3L7uM+RlNwhB698Wzg7cDJXistHpEJ6hA5l
jJhXKxF2Ro5og0qwLZOtk348Sz6lwLTKph0qYdOZV8kWtCGvNew3pweQNn890X5Lvayctfi37lmr
nTnwBY1g9vqvmG3RN9cyR+zHlOnpfee/e0buk4Azc+2tauuIptVKRM26hiRpgsuAFSw1Gujz2mq9
C+PxmCmEpWqinfSCcIyKITIht4ASoO2L8TPFlvfiCD0jS4hHDSx4gU8PnINC03d8DBzVFjtliw8Z
EYAAEiWKg1MzFaQ8CUZ7l0DTua6b0q6lNmr+xM6PGPuGB9vyZFob09mIXCjgIyxkHbzCZkT9b17z
sUkFvy/TMOEfiz7zrKZaFgQ+F7IL7WPcrfe+LVXwkcp7MGouxVqIkUgWnjW6nH3xe+m/DpI17iQ+
Vn8m2uvp9pS0vJxXfKC7jZtemQ5DOSQAATiPyKqxEFxSgSoyrozc9N+qzIYQwBj/OAcUJEL/HXFr
toMQV33O9VaJzFVNoG7GMAGIcYZj468J/kgFJ0sEYgWdgQp+2fIAP2ilVVHfRwdMO3PEKgvKvYwc
0RTrZF7g+/pQEQW0g/7ARRyeV2zpquwnPTu75vHhbpkAXSjc6hpvcGBy7PSv51mCPSaoE3MajbYp
R8Hgbm9xKvQs8dxV6qCtKgIn5VJVKGS9Yc/9ayugjCHo1EdmMkMKEE174ZUFpXRekn7MnrCxGVmo
d5QYS8bBZrlkrcent1rpRTnfANeF04g32SMfCHyaCuuf/fTou+/n8luhIbksmiUE34ZvX5weBxo7
cmvJSr/kIeIxTHSPWv+GkS0V3vyraB4RVZj8tuv5CKQloc5A4doLmljAk3SL/aIr6LK8qOomZPol
VRjhhwf87mkj4h7tW0gcP2WMF9qHaERsW+Axm4BZdYyy8YGgQwkiKkIwP4SqrhmWtA2uKtGoPPHo
kkB0+E2j+1c4B79+khs0WRy0NJs0eXXTmLraW4m2p58dC4ZwjQvr1evkrgtstPjcahYKJOtM2fFA
0snK0aLbov6J90C6hptytx6xKbYG+IaDtbVrwLA+CGBAIPkGXUoDQbSdIxzN3aCycdh2VG3U7mzU
Zv3stdBQdubzHQFXIJCqMdRkeNaXBaVGaLzdnnvIiosCSxNr7ah72BQuwFhdRDXojw0sV0Cm1okW
ZFORr30R4A5ZHZyTb/vzziKhN+Go0Xu+Fm0Q/NyeeQKb39SnPlPQjIwd/8JyDyQEGBRf+DLhHg46
sM1vLGKolfuqdJq7XCgYoygmpF6T/rt8rnk7xmS0dLgAC12Wh29B7moIvTe3M3muAhLmV7WxDOuH
MGqEl0lj3jddZFAl54RuiqjRhTLd/Zvyh1OahZXJiBKcqu5S4fsccpn8k1QLV4DO/kZ2YxJ7gUsO
mYOK+D0zx+Q0Ux09CUziuLk+mEG2SJuSGwKxWOhkSiRhjy5L6V8dBZnHH8KbRY7LGPRilETiSs4J
4v8N8XG+RI1eU11e40/rwMjc+pjzsE0JP3gqqEBVyFavSxNauuSJCmOvjNHii4t3MYt89JM1Gq/o
0JTop7IhDKLI4wBRBxj8NJ5ApvL8214rkw5qWiLw1hinA3Dryl/XQBi2d9dBGo3PetK7mr+jVtws
dZfKnaCefKDm1pWI/0qshgJS6xe+K6KbaMSfmuMSqfqjdOMYQ3ETJ4x4tPafrxDKyRycmcFfNGET
J8gPepNjbyq6jfufyX2Sn/BWQs+jZ2MQkVVf9dq05w+0ogu9FhNh2vLzoHlK0T8nDaj3H4tnYe3+
a69LMJnugEqLIlV5jAwmAZbzAoJS/GuyPgC7hOsvC3tJt+TTpDt5G288cOJTOTwHy833dbK5nnWm
MsyyXAikSQOYpt4F6xJ+sNwF297Y1aAtBQ6QdspnCDmCRKfww/98NJiuletPDTRRVo9gimaigZxX
2lyDpnGkgFL0v85TzYdYd54JMLu1Z593V7v5o2I/D3ZGU2NwNPEOOcCd/J+HbqY5OL/1a5rXaWnJ
0jDk/3OApu7NXJR60f0K50/XFegtwpDQasN2chcMLWBNHQHwiIqbQBAv5b3m/ZoQKYenAtSjfila
aF97f+KdTHjP8qAx9j76OZWP154CQ05YOKZnOWF8yVTAEazuRmRaszAofW2Xv9ZipTE/ro/fz4Ub
p3KtRlGQsl7vNJwmj7PNzAJK72m7uHTYSOuZsCJlS6T+r8YSmHkawixgTTmmpGJhhWsL86g7ajaU
2TtuPIDWpDbkjAA/8zykyoakBtHrpmEcdiowg4ShVk2KWlM86Sq5caXSLo11163PCE3jGB5gSSuy
Jf1tOueyqrQhzKY6rXgMkvylgNe6vgFWabPTvCzHY6hkdnwSWmFkeHgtZdMmgJGua6a1wBNY9BV/
0utHh/xfQy2A8dMs5JBKdffLNsFIKSijR8lpMi3+MUFoF/9pegAj7POKgmretz2ycjSz676W0+fJ
JW9rJW+9NyBkMtDkjH27uOYZpVLTsN9ZWktEV3hEo27/CI1RWJivi10z/1TPUFBQ1bNefkWgTmJw
wDCPwpPr75KXFYIvkuG5vsL/g2mtn6iNtax/5PuMvGBHmL5A5boemEAyetWaENBz4s30YsX4UXZC
p9q0nFHUqVxUuPymjmuIyH4ysl2obUzOeD/RMPIV/STuyyfaecJwwKeycut+Rcht7eWi4zDkPuNU
rtFvS+40ui5WrkV57JbumJL6SsGmRdYAuzZJgC8yLvFDj3CFCH49ckEmDMLjFOP1DZmxbSkP29pt
7tXaMl/BosaBrHwR9y/OipDJ/UGHMw8QCB+Ip8TjJS0XZDetljAWJswIaBUfyHhZsr+e82dxZ9sl
16n/IyYU35cHDcnBu3NHEi0PCYN9y/t7JKtMfLGiadNSpKVu++w5sJENZcTQOza27Vt9R2maAabf
/kdm61tx8utUb+QkgyDHX0M95GkXUek+Auc9r0zw21fc8qMIRF2/ys9toD5FiCLj7LbEEUUOOB05
S0Tm52JSnwsDflaE3UrjBJz4YoLdvg57mZAuC9RGsenCwCtc9+N0JqCnLwUXp8mlZxddSHyeqJwo
+Bht1JLL8u0Tbfb2AEmAkpNzQF8TU6+DthIF5rgmhjU9SVbBzn2nFW/NXKCLp7nJ3YgD0jUo1xEs
dNVlT13H/itX1wlroe1xznsG9f3DgdVRiocyFK5TGEi9FUgTIvS9wLO5ys1Di1ij8A3Q627HORTK
uejEXz7Qgbn5tfQFVbpTmpD3RJkyg2iX2kD4I1AYsa0LusyvXLoSgeLtj4bQ7DDh1k6Ckdrz9xtj
8Fz0x+c66Zm1H0gE9vPj7wQ8vsVfCNORYIcZ6oJwnlVJcNVzyp/yfwb8cbKmNnKJXt0U6YaV1zKu
XePaXatIpOPwuyEuKuSRBnDDBsEdtEGv8qpIxbinN0fU/IlDd42PEfIEsDXXOPh+Yu9zODyKNPrR
MXKOgrRohRHi9lQHdo6fZifNZgzMITWrJrQOv28nfaa+5yxZYzdF+Svuz14PRFMlULDV/TEqkYh2
c5gH6G8CTv6B/e/PLGTRp53bmqBPT0vFp+WXJpxGEwAIJt8uL3xgymElaiQ8eq0XnqekzaamPSIU
Tq9StY2rMIlW1/TvKLjfRuh5o047XeeJuAO66vjRi/W5A3+L6v4ej2WbqAPeC8fGO0IwEu4p6cso
sJLZXhcUKPGlskF2GlLY7xgovoXaLcRhb+oB61yhi5gEweBhCRpLfNmk2vIUSQzTZUsdlZC7rhEK
HC8eono2tVRWsguWkhCWN7yFrFtMRVE1xV2SfUfzJqqzzhf16R4zRGmAaPJ5XOanrzrYk7tn2oDG
qYHqmktRWEimnmQ8YVEYshaWvl4zBoNULL4fqLFBreY6/sHWBI6BUGKWbaAiR2LawEXRgFNTHuX+
tbH1s4J99H5O1xI0pT9Z/ClI5qyEHocaJQH581EoLXQB2adn2sIdvgB/sdjE+p++tfpL3uXT+lTT
UwXlh+Bq0t5sP6RWvq+XtkkbZL3IUfH4RAF2Cc89JGgMORBWmN/X9hFoqDsbq6lVpXSk+uM40/bS
gwscU/MjDVqyQZ7r7SCAZe4jvOuCUjKeADdCdzGRfNr2HDlQuBLjo0TDHdWcDhBUhVkzitisMg7Y
ae2TtqCzKSsMLiwj61BCm4oAxZ6Pd2puicTLVyXb6Oz2Nj9ouPZgr8JlZQEJEXdGR2Eu20Hyaqoj
ubcEZB1EtRnev4q0Hsb53490FMwrDeZXfqvqwcAqLv98Mebjvq6QqAUDAVMmzh651aIumaJ6bbF7
Y2zr3p9VnDAxeDCGix2PhZEVIf1Yg6ycj8nPcKy/ZJYbShyvkUI3d1iMQNtH9whOAAYVRyjKrmKL
cimw1rffvebcncYW2FVMHj6DKFqZx6rZ8TgX2VkJw/1SB9hpRyspon+IaoBzWNdWwJtvQKXbuMk/
/5/XZHyK7X7H9QXc39CbBkKr5WTvXiBOPxCIAcIlmJbBOjs1eVR6T0HmvEm0C7YMs+dFDTCIDZ18
XSvww0Ld/o+Pl5IaRj7ANi6vsQpqW8tc2ekZ+17nRiqsochYcceZs+CnBcwXfdaq4gqZaGvuSu6n
R48UVaJcBcodCujrkgubZHr+hINFGcgPU4T+7IPz/63MqN3kxVC6Y7WkzuCbUC+VpBll6cWIUzWM
7ROPauizVaQK+3/9CymFVW0VKhDtiGEfVFaPFc8hO3CvzqQnh1SUqtZv26SAZvdYJJh1RQnkIIgY
OgFyBByzldMA+v+M9zSKW9TNfhE2gsdqy3uA2dfA7+Evf7eFfgfn/gIoF64JuL2PHAZDAhy5zR3o
axyWa7jxVK+aeAlSIVYvd4qg0dZ15quUGlRALjvTaTVpJD2VsYPTpTC0Mtsqc/lh/pL+in7/GUv2
v7yBG1Hxd+ejaJnTEiuL8I3b6otfmLsqFrslfyWhjascSZaczos28ksa/Ke+UpXGY6RPBdIvRIWG
cA7ixTGpIn10d8u9goJfSbT6akjfzlw0A6d634QIvfw2zdtJQGNlLDoHD13u9TFVIxgut+k5ZqcT
3PvifksMS7+9eqzoKKwBeqMsEbtkU8snqdt8VSqFAodVxkX0oxp7qW6Nz70T0PDpbGbEUsyCIK+0
O4YKkAIIRWIfccxCffSx+COa52BuIkY00mlFNKyOZeOacZBMU1H02dGKtFhgpb/zk5vvI9fUItNX
SHw2Pu04tbp7/eE/eqQxuf+uVIAzQI3bmqSWmwESa2gymP2wYNt7Ol9RsGvtszXNvD+K8TxrMyR9
/KxgkFSOjtC/xWgL57l0qOSghMO1LDBENmO+Lz/X4VRocJ/eZFHyw47Xjq1jPH47ZUQNvFEUqdGW
M8RTacPFdV9Fh7BXEbgeBGgXzQCisd6EXrExSAgQ6SMvA/OLxwwPXPWzrYeloNMuITXiLt1SZc4w
wgnDcUEIga1SrAC4hlUrbQYqXdOqpwHMebWCC0qWhUb752X3x+2ieS/vaj8RZcPzJfmyGE70J+xv
QPnet5J7gnUHCpsKyA5OAbA34eF+KsaeSxjmguiBKrV5ODgy8z/YPs2GRjJt1/ppu9VHFg7lq4q0
HFQNap9OOIYIZCIXPGxqSXUsmBQpAwfjnLZxUxkUqwCN94rhAsMVAevUZ5JLiO8xGaMjMu/t+UL8
RcmCcFYn0oH1mooVAzTn8g9YKF1M+72VlVp2CPOL9N9bAiBuFFTiMRz1HXSVOTnPLX4KSQVsx9oj
TqPueigjYrYHQMy03Zshq1pFyF1KXk9MIYxvwGSm4FEc9iXbDq8Blc0LSl+VwOXFUbgSngQ5hctF
8UfGhuFEvbYCoeacpDB6XoIU0ObHc+KZQljHh2YF/MnNSZhu4xKS6cCdQB3vO2RpA7Jp/M4sGuL8
vRhKykJU/4Aq025az30HJef6RQ640LIk5LfvLmBy8nn5nHLYiEsl2APAAHDkeSjvBBHqgDAicoPB
QKZMGwVcMMZUdZgHylImdN3NxmgdoP/vKuyzdHBE01cdkdRFKQM7Ob98oHCdvvQUq5PAFHSpPm1V
WbyDoEENz5zkCBftiDG84axGWm7r2tUwXZhi4Li0X++CtEzlqBbgPAyrdWodQFcEQQhXRWaofbqX
tZa2Iqnk9mMRTjT/Ri2oSvkZb+CbWP4O3mQq1AF/W4aS+ArdRNu8nTWiSZGRZ80yiT5/86X7/q3z
cne/3/7IYv4uY+sxDlQtVff4XWvvmeS2kI5yelcMGpJPP1Yuo8BbWyjiI0CZXUDsAXKSlpPRYVCK
j+dB2m3T+vRdv5I3GwovtrUwz4oQDoTD1BiACXst+/vz5mdivxytQVKtonMKdrYxgDG3R8I4/7Aq
XY54VSq6rcEm42yOfwXS+JMboEvy/xx1iO5BW2EJygqpWcYHw1UsSTkGdeIp0nllixPmO+GrGEQq
r/nqnhM+YvnU/vpeRYZ3PJgwSTXEY+PypULAsQA4jZVsmwbuMHEdVmZrAY8O9LYpFQsfIOfldJRK
r+Pnjo0deLOvMWBbybkbBEmMYTo3bp+K9D/Xo4oL/6tFEoaAOSgUcxscNxE4wdGQnp4NSI6EeYi/
NhXdtsc8Qo5neniyPE17gzjF+ORxuSL6EmXAEdiBG042MfPysTpJ+K1anZlJTSJyRjm8SN5SG6HP
ShTpDTH7fk1Z7xE74YuWAtOL6LKZpSlAc7GPJ9kGwROrwwMgToJx7xixlFkkAyW6DBQ5MCMmh6li
OP+FcgBW+8qRBR694jKZ3V6j0hZAAIDGZGCNQzMCjkO1tq2t5Df4erJZsML2lzQh7O5sEyDToqLn
q8laMYqHNH+ZA9u2Z/toYIFb3Oj5ECQm+OniqXL3/JMC+laRGKEZ9XWUKqcf/oYJajhIalt+M/69
PnwNW+rlmhjgbk209mkr5SHBpyP+hKsACi6+MbV6Vj+HXsAXKZglDu3IrXP4mIGOSrC4IaiPUCX4
TBohCycG1Z4LN4g36U7MnOeHioT1001zPlLE04oGy9+mPuWC77ZJuLtTXJMnkpkyKvCbCehJRxG9
JLvMEzDnKHFjp1B/DWWw0gyC39nvnH7RumR5kROfHHdkXXlyXEkOuZDO6ubWIBwNSkVLIxFsCrw1
dawAYHNMUm0mlHJJLqm5RZwo5Kwr0mxL+zea1QWpsHQFOwJZDL59/0Hbcv+4pHwYZBpKlss13Mgs
Jd0UOnEc/bTA8HlHJt6kwFEmQ7DwZBs8xr9lIlgLfyvGfZAN+Xs7gIj/eB1gOWABGUB5lyHqnaG/
Ln4h6tn2TWF6sjUy9nUg8VH1Xb3fjXbK+Fn67aOPbb5je3ie8YSEHmIGHznIUhgdOVrq+zootc5p
sNjA1n1TaA4h9Z89XoHPLBqY+UlXNUcbgw25T69t+4L64b1lBN6kw9eCweT4EODLTU1++aeYVWxA
51PYeHQVmUr5+4ATQLX1jP3qV4mTWSMTPHcSVKPmQfWHr9bz+ft8L689y7ZzIBko9UA4gxdHKasU
1iqX8S8AyUa4tUxEeIj/zSRJVz+PrkjX0cIIuFaSxWoreVtAjkTjKUxBoa7kQxQ4vuiODJuhrU7K
geV7Lh3Qn8SluOtmE2jKluMtIBbVNEQZ7wv+VZmXINmRtJLxkzdTthjn5aRmN0iR4LgVLNW8OfBO
RycZWSLrqM1YfBHUYf1rgn/wcr0Fmx+ehDYtKesrJ4pIJZWjO9JXRsA7YRA+Ozj4HuIjV+y7zU46
bP7TYjfrQNHCwx4uYwnyc0KTS28e1nseagMGqttx8UQDLcnkGHmrMN3ykuQG33BFqb+BRKF+MTat
I1qhjf7Jzau+9JuLGtZBhvKpo3thxYdwwdWbfhtR5d+PVW0LxbuTyu4Nn6B0YzDBJe4g9EIfuXAo
hf54H7losBBzhiOpgHEzqroBBAo/EjqAL4x4+AKpap6K2ow9NhMsdx6LTyytS2fjftXMOQsNpGsD
w6UhKngoPuubNTQnBEj01nnA/Y2bV9xnP4f1gKf/aRX4nre6jnHStSfXh1F3eaqWUpPEdfYgXgKy
96V/7JBrXUBzqxziPxNJM0HHjUwOzSWq3jx1P1WxQZ7Fkb8DZzXm8QXOGYxPHV20DkJS4NJuMrfz
UNm0OgFvgUAKXeRQZAAi9Ascg2lSy6BQNonWyOk52yss3JybvFTF7TckAjVDU09qHrKfHxdaZZZc
5oJBdhj+6gX8Eu/P988jIaNtNYxqkGb16WtqFLjrUULSQ/UMTUaAoTAps/RmI3s3YjVA4JcISCL4
gUBOfYti0cMVIgZrHReqO8a4jUuyFZ+28yr7NF3B2ORMAj12dV2fg9ZjcDVyL29OM4Jk3631yaNI
r/puAEuGW983a9ze7EHLkytC40R4w9rbTvKxxP6LqVz3r9OK1I0hPQg7r4kS8AHSsfy3/tYvjIm/
iG+1ohzzsfmwsZ62rMiWL81wpxotlYtRkiZN9COaQuz28MPTPr/qGU9pLhKPDzimX025QYeFjxTy
xZqGWuQgnXODpk6DgXcSZ8dxpvPzTFaMm1AefyZU2ZHNuQIt09RlYro7uC+NnoJ4sq7S3j+fnqPJ
7u4PkTaKipKQnCyTI6cYipYxe2VYRIT7Ykz2gXEnyDwy6VgQT1RDJMWco7QHS9SWM/YBQo+uVq99
SM/AX8lITRj2U3v2LPzTSKl/hVN9zhqH1h0/FC2V8OXBC9RexI+gC2WZyjCt9noCgTLEU5UIQpQZ
ew5h2KcP+fXLBbHZjOGD/r7f96OgyUMwZ6fOEjOpZSlE6DqgXAkCBu2riZMGP2pOWxlhnlBs6mNP
6evWSaSjij7uM9NUYkeucmnjFPGgVwcruxvQAplHiyRn/5gDwtZ035GEz7Wk2l8YDDEvCx7Hqlf0
rmWdW0Ru1jVDmlh33sELYYg9bHSynulaL5CjCmllplyqLwzDyKZiAVZHS6HVP11iIz8j/SjJHSn+
UN0gBIwnwVO0y7xExbNtIW6nrqZVo45zgwCanRHFJmN0E1gE8oCGo9/bdBUmAsRR3UwBE3/wr5Gr
O0FIAwvdoJfrQlrHBurc9AVt1U2yO19Vk/JI9tX1K0woi+jAX4Kn9LQUfFFZ1ZvoGvOd7YmbB3HB
YTVbOOVIfsAbxUHMpRwJH3UMP4iwqsTurTQkLqAsmgubXAiJWDyhDD4LXL/SZrqMdyx/IDWbdexi
RJaVhgyzM+gq6fOIWpnXl0M/v5INbbx0OhZWX5sLpVbzQc5mgrrMR4KLN+n7IFq2yrDgNGK1xmSy
TJ6DQqLZEQnqyCJ9+xLsXyKYF3a/wvAlMmYLmCF90Wg1PRkQu7YABZGY4ha5pzgFvxM9R936AXF9
96tqHgNnhEUvg9CgrfUmKZz5H5KeiJKpQGZi44iEph782m5bI7HflUcYR/D9xVuq6vyNP1s7dnMS
r1GVcQCHVKQyApeQlLNeuafuJnMesMRCekm0jUjCv9FyEFZ7qEYssIkF4NP6P+1DlQYgC86MjRLI
dWpBL5m3p2fVxXQ3RCOUqdXAfy20XRRv52bBBtMt7FWQzPIXLYiLSFJWJ3rtELc8L3P1EjaU/hSW
7WDM6uur3fLu/8+BRZtIcOGUlA9FLTkg8koyjJYQwkSEtqp9BXip0a9uxyj5lHDjIhdcJ7Gltbs5
p4CHIhkXFpTcMNAuk2HNEOS5Dnz3SgGYXzWeWasxbkmmdh/cIgVPGg1Y89gnQbOsqjQZPyK5LKiS
OYyntWr23bJGYk0KBIanp8D9HRCkbFmoOhPAw+w85SXYdLjBNlsLfX+Zzf7g6tqUEDDVXv2wmGB2
y3mcDtWzym/uGVGzM+e9thIqaEgUE/hXcTwvEw6MJpDrlELJ8g2xCTuIqgjzEp8HmU2/6Ei+beLp
zpX40fogkUFpo6W5enkc8IOY9ag9AG2agkZ0RoX0xcZTuAAsElzQC4lBSW3rQYonOLdydMGydPZz
NbwbiY9pNl4gThw00U2bz5k6JJ5rf9ZNkLxakT3TVk/nCmGx67boSVEwVPQ0wt6hVPb0AtfxRnHl
rdTdt51n6WgRnakEPdi5cWe7TsIcEYduf6nZ5BcsGXvoRBN9a0JKhF6Po7bl9DAIEefoicFRcQgy
VTJY9eT7egyuptQjHy2yZkqNvTO7Zqtt5aSxVAhlH2jg91FqtwUksWy6Rk2DbsxeFArZbi9ZQnzK
UL1jo9ER3zwHNdWvRQmdkMjGGAFWnutKuCp4BVmlno3XLfOECR4A9hhGR/GTrZbPYk6GUHrUF5hF
t3uNQdg5paerwd9g2N+y335K7BJyFINNblY0Ewsk3eCDaMTrhkRH2krocaqsOECvwiKHXiWdXYqi
WbCUZVWvX+ZbYrLEx68jYyRGuZzF0FxfT/ZEA4Q8LdioHhm7BXYBDhYPPfedfZWA478RYEtoyY7K
TlscCBet4ojV2YMRifS4PqUb0053+Xm1f9jeon8d1KdxwodF/xm7T02QpUhWJmRWlvkywrG2buO/
OEkAuvs0X5ns/ElYypPEvi3YSz8GeJNMcwFpE6hScm4ADy6WRSJ0PB7gKuCEgK3GNosR6SnNyl70
vbZV23mgVd984mWfKwlnlpw4BFSmVldLiESwItKJtxKhL6Nj2KR24hgaHVDsPOXqQJSe5XfhPYct
7axiLhA0t4P7Gz+wHcrl/qbxCmEfni9aDvsE760XD+6dpiC0R8KYB2KUmkUzi0Bte9sIXRRclCHe
xGTS4JzPeC+oBmI1POrhxq+ZlTwLxZqV+3IOlsviblPryZkeX4EPSOhTflM+QFCEDHq/WRRAdHKx
U/EZJKy7B1mjMF8CB8KkvFtN56tAKOvo4tDpqNm1d+iKFmOZHuswx+zBw7Lsx5Z/gFLZ1W+ooS/T
eHxmOOXkwF2N99eV8RdOlPr35b2v2Jdsizcq8j7eoFs/I9oHP36sNWkukTmfMe84pms+eUqQEvXF
lPZ426m0ZpL34doViO7iKydgJ+u8GOvECeEzYxWaLVV3f0yJA+knf5OJcDc+vkH1uDAf+4A65G/T
2GHFLNzUVWc8KVV5mPYzOZ5D9m224NFf5f2eGDJzUXTpCPcKWn/WUwoN1rzMYrQLK/l7IqcmMw7e
VYR43Z7o6Uj54t7F8RDabsFNwtyHcqDuH9zC0NiPTWQKKsMXH0Vtd6DPB4owoNi+8HD2KxX6SY3m
FHy0Mz9umx8yxm98a2vcZbEGcZcTlFUgM/upH5Og+Mu1Lhs923qApQqfSq3ptS8DAeLGO6kvHrjJ
+nIPxWAcfXghDBE0WjPuhSJg6qn6duSmy2GtvAs4wsDlXKsQN1KDKiEtxLskhOE/qN+J6AzKhodo
SHHk6YVNJZLyreKb0184YTqA/9yHbq6qzRCg+boa/+wNr6E7B2/qts/nfQkBkgpwjTSCuXW287Lb
gRXvEwDFAuIoK4bxUF+aTiN6/A4CFjXjxyt+b+AOmVzzzNMdEME7537S+tNGrfZHOWDzTljDyWA7
Zokn4lPibffLknwNjykqjmOoPCBg5r8iyGPUhaHUBehYtSQvQdbFYSBJhPrclcQJaF33vA+2BpLR
6gbyMYuyiVC00bs3D7RQz6iWeqiSxr/3PK7mtvLfsNTpYeZpH38HJrpC1Lv1NibuaFmO4E4zj0Ue
hSImMub2CNY1dAZCCU6vLeHumF+B8X0jqrU8E0aRuJE8AnQQ0I49ltoIAPkfHV9sBJrl0wNB8JXm
tEpguukgUQGpQuNJjRMGmCNhvqkDKALeJchzWBKsqBJxadYSIABxOEh92dQKyOHZphQfwZlXjVde
laJrO7YH2OyHKwHsaFxgqZChYBl5lAaw5SML2lcTSfqYnnnvDZe0nrLPUre6ZupkXbCT7wH8e3jH
WwrSnDcrSDxoaRQ6x+nXVGurOFMVIUFjnk/qyQk5jfwJh8wuZpegxh7Qa5ORvYyK3cb3W/nfhsR7
X1TcEU9fvqT7tUJ3WVQkQHhtdvXdAtjEKfwIxET2IZ64d330Eq22otf89BYZUfegyLsptCLkJ6qW
9fMYhTkIicsx9lmpflv02pamCJN3m9k4Bx5yYXNhcNJ46BjC7fWlCqjhDQ24hnrv/NuxRUbgcpUW
anh6x5TBls+6Jn3TU0JFimuCte2mQkkY6+YCGSXNHLOxlYmnd7j/eaLs/9NZKRrLAk/UFeEF1XdU
ZjZz8+KpqseoLtnof9nE1IFRNxtPtJqubzc0d1CzE873PqUXg9cc62jcB+Ul2jGtn1lSFVrfEhxs
1iLB/671lzW+WRECKrg2Se6aU1csbwVl6re65CfSiHwkJXcY0ipmgGXH86q9Y1iSkw97geJfAnM1
poFOlAyzmZ31KmwkOug+7NtcTfGca/oAhmKwakJ65PSvYaX/3gfA8rX0+63bUjs9Wb4HuivAjQMR
HrF/G9qQDFAaTzuJ2Aib/nAgQP4gLLZVethsm93BBSCwu9LWELPVAe4mX4SyY2p7glAlEGiToPM7
leDCmFUOAE+BESG+tlHFZXazHdNjNAV+ELN42SjuaNlGo5YoUaUg5Kjxmv2Y/NH/0CvOvQNQRpEF
PbqckGY1p/tUayauv19GlxLzhPX2P1KWxlmlYA/PAb5dWsT4/KEzQabyuvxrTjRLlAaeBB+o/O43
CTGbpkzI9L+odkU+p6rOeATPLWI0b1dh3wNdPgKU1PlYTvlt9Mxy7ZBRB2nlR9Jzlif27+JYaNNt
Q7w1wgfwagrs+0U5kkNzvlpgVmGg0IS51d079rtnTV+zVq6U+ADeKrCfa5fFMqn+V1r5/R2st1Zv
uwGC3gKj78PLSuvewK4ElXFoLMSDwcVHs92EDJwigdpOVsJjmYv0UXGGXbJlcOOq9p4Gy5ceCojX
6gpQKYxso3dPmePPXGQR69nNU3X4iKIjrlOUVL7INx6AGOANsqjWFZzgkayMSmO3i4no869Nsbbo
WzpeRJoZ2UediZr7ca51X1mLEZNM5mV9qqLlU87+XdZSWXlqUz5ZM8JbnHwvqDi2j+5AWFlqqrwq
gUBH4JClTCQVWS/mZI1XNT2CKKGFKDIlnw362UhXJL/AOLC59WkD7iWqMfPxrAaK0yQWFIdH3TZE
H0c0XbEreUzgYx4zyA4WPEyhxc5GJlQEqli4iItSdDNHi+J3r3x+wu0J/qH0NZcNDR1+1sErBw7F
ta+189HXglWS2ZOsFF0OnjY/vwCAuA11HLjiHiTOeT4bcEl6UJMLfodemI5et3I3uTnUZ4tsnPwO
ShrdfH19HNQX/gD9E2E9ggQif5lEllH9l80RYruhQ8JB2DyP+Tnurr+yiznhy0ntUZMBbXNYvoxq
iBrk8nUgrJm1CKCOG8EVJpuCd4O7MLuw1kuxgvGxTHKbfofwvmmVadpxCVe7q2+MZr3zR8VqdPnH
QgC62rbFvzCJM+2OWjd6u6SJSb64w90ZJyGaP5SY1TOM1z4Wcp9P/0RPttX6BELET7J/Qe1ZAOPX
5FYjb21G3+KPZwTzKlkY1o/IIm7gFTe3hCMQiH3hrqxY2DR6qIPqrqWrqrmx83f7t8zhNGPRty4N
GGUlc7okoJxu7Fdj/ahRGVvKVVLEJn+7+oifkJIDXnA4iwQAF/AK/ujp40IHKSmUX9eHlqR6JhOA
1YQPj0HH5qjBFfx0HOy6MSaACxTF1tp2fb8Lt8R6z3p8DyzDkZ0xOUAThJjtP8kBcKXcY0SO8DGs
UqXJMghMsH8GeOruwGgT69DQHaBHpIXpgv+ETtZObptD+m8wsqfeCRj9J2rmn/IaXaecwItN4T+q
8SCWKxmB6P50xpp7uQqFajVz8gfzU9bX2yYZN4I2k2sQcGCFONfvdFagUcn8RDeN5Bj45oCiYxY4
HCEChPJlIonteMaB4+q+yrJ/L23LmzFO4u9pAsECw1+DF1KRS2thSkzVLoMkP280A48zdUKFVUSQ
WZD7A/Tj0tZ4T1opGwn/dhX0+F4LJcqKw3We3M6p1s5wxQpi2Z2COkihtFJIziAK7IF1oz4wFl6a
FGnDYB/oqy6GF2yvuV0mc0wBgv90XsR8zri5eo5OrkA5x6WtwB/StxwXkm2FzWK5ElsviNkJKrWD
jIaHTPYiKOHf0hImLxbN3i4MJYA85salNvyHiDnc3DaH6MNYSnyMcsXsDc2u9ofN2CHA4czarcHm
hSwgxKZA3r/j+7l+5mV0Mlbt1X2hfalSJ9pqeV4kgrmMbiiY+m0HGLGITjr8+W4uZj9sp2h1GBnZ
OfMTPk7EL4ZB+jZAu/kRJk46gbTj3y0sX2JmIPIFjCf7b+AlC3AZarfTghGmIJw6JMNHCxErLqi/
V+YuHA1KmHqsfazjpul7DIT8VxQ1ER6qiyRyehR3nSyDWzfm1aesjpJkK68AgnA9+Czhb6Fvr4vx
NTSidG+QQDRX9pxafrntm/gs7NWs1uHVlKvSUieERkHaUrQ00omeUX8X6xrAK7nrr0I69inW8nyb
CdHjZxFfve8VnNb3F1ZAcxcFSMwin/147F4FtNdxsWUPPd0pGvSazNkZXDvH45Y4LE3LBnttnN/x
bb1LgjnH+kNyC/mHUtXqdkORubvb0ONUaCqCo667OmUFLw23yWaVDbx6h2Q2pZd+JU3gAnhE5L9o
M0Z9K6wtOUU/3LU5NT6WPIveTy6Z1MmXVVgdXlfUE9MlgGEtQOR1wrK8/zsMY3/OZ0zdbNW6lJR9
CmVIDnO+HM8+R965E9K+9U952JstD2G4Zqx+acVd0rhJ8H9hFAJ3AY50/QtkuabtOcrDGYEOZhlU
4ODIerxV8cuMYCXC6x0m81z1oie360MQ9q52NqKJSnhI8ScLUgBfe3rXDfG4elWCFsmPn8/8m4x5
NX4LKomzXDcM2aQeLb00diVefT6Sm9I9nVh3Ccdq+VHoX58Aa4IxAzeQupTwZPHtKzgP9BnkqJfZ
xMRKgxujI5j2N5A2CvHTPaPRBYZrTv1xzz39iWprfQmxYtZhIaqmOvlnHbMsmmsLI2ZJkVZKHCnl
r1Z5azQ+Ow7dBsm0xONGCvYXtb21/jgWNE7xLknsGT28xQ5+yX18Dto7XdYkFP8smUFRe5eBlN8Q
7oRtLVpfCsHawzurPmbDCBNWPGCP4mZ4msxHZUqSqwbS3yUR0lfze2cX0hjNvyQ8c3vwR7Jdwtcy
m4tk1S1/AaOgfoPqgdnOTLI/6B6Pg//IcJOcP+8LNpvONDui0BYohTiqp2ZengFZMpA1tsyx6sLY
r2ykUjoQaWXG9LZ+nTdls2TaD6RjosdgzZTYymF2pyofB20y9jSP1HtUXww5PfFPFi+bVnFfwhrR
om+MAIIk295+GJ8X8f6bW7S3HHoElqRWntEDQcLHl4IAnnQTTbvXEgXbPiDx092gy0vhQdGSMNcT
umnM2NLfCppX/Bz4DxYFy5bAGORt2UVGtGnms+e5dk8K22EZi9bnAyZexlaC1RwsQ/ngv7Py6Gbk
6VJgDn1KzD03iUfvnvFR5NRow2TWSNEM0FoXsJNWleKaXOF6JLGfzcLT20sY7utdWUbTE2aX/G4G
vYRJU7ELDRjONuW/CJ/kWZLgnFe4AlnhPN7Uf7C4zi9k4YiLC3jlda5nakswiz5Sv/buV6EikOsp
dpmQqvrn5x+7999BOR3TVDB35i70evqFENEoOqrINHvIrd3JhN817JuO0+NjIPqLVoX8bAVsTKeO
jPc/HgwHr+81rrsopr4v92kllB6m7wFFvnvCZOM/8RSrK9aVg63jgFoA7/rzpEWk63nUeWjLkga+
3qbW5v+/hJ/w4CUZJ/xvN031A583hDVqh9J+Ec4hOJie3gbVKkUiE8uAF+S8uPToWyyPfusYyAhj
1+K7HopwTol+JbIzRln6DcoX1kSl/ojsDP3hnTjy251TNQHvumhC2a0SqxMgXjeozFrnWgwt8NXA
McsjVk7W86weKFyXNgMvchTlzxtCNksKxqKXXJq+/8fZQm1DhF1aC+n5ADfkwNRl+avzffwpF5AO
SaohlbPoeAtXvX4QiaabKqcg9BQltyi0xt5QW+9UiHmL+Xfk5cOVNFz2JSGpmDlsgNVhnygP8C+e
vhFLU0JLneaLwDmolUvarSJ8VnAQHbTGpO6WT4xiqucEwcbeLigABcNaCU1IVbNjlQbps8lw2o7i
RThEZcnF72x/22015zRacW1Sr2f0q/T0kCzpC3LPAhE7Jl4KGZcO9IDSr6r0b4O59mTcro5pHpcS
PgGBnyZimjYL86nXBnHRdgpKDONaSPUdC0T3iDDKYfyZRWmnHReqmqs1EAA2lmxBJfi4x8AaV7CN
2dpfusnpH0YvvNL/Z1vxc8AHhemYqiTBZctucLCLfDncEf6DDd425lwjoRzjTRGEcNoTEISDePub
L9eZcLrIhfuF1XlkD3HeZ1sXSOTVL8+qhsC5IHP/kvjkgJ8oLW+pggS6MiOoGKv4fd1eoSwzvJhY
1mL4LsiKYvxDWPpvHqL0ughCiJB3nL/yYnbDuaZYuyJudZt2XIoFskLR5RoMIxHKUJDSe7jP6rXu
RgVQO4DDinwqvaAEEjVVyEivepwXSr9rRwp8b5fUmUOk7UegvDZU55hUDnG8EJKbSlynEsPom4sG
vBdJnNbOhMu8WPfUU7XBD2eKdObVs1chivvAE+MQWNwrNKjdzFe0zZ3OlLV/GElxnfbPlw4OhN5w
/E+3+nsg9ojnslBebud77YIBgGZR6p3VOSOQSx3cg1LC34ZK2EG6p/l+y8FHruKvRpDMkQNcN6ve
ydXBlal2v5mMBt3D+WWATMoz9vdmKdzHfld7c7wre3EJa8EOivGLLM6rzj5uc2rBOHnpltVWDyfr
3gs8rWp+qsK8+WxhnL8MztW8z5/D6b3S86rge+ZObxFtDp9FucUUxThhd6oaHDlmXxOVZUqHUXpH
gpSTGFYdUdkw/YgwfY7rue69/Rp0o8aS1E4ehJcrPdlCsYc5rMioGg/kqpdMPPhsQ0NcB+UKji77
UCzW6gXg9ESTvXPFKiXCN3v5vFdzxvUJI9B61yogbJQp/acVdbqnYUaYr3pdI3yjJaRAZbPqzAnS
IqbzEO2RD7sj4fpefltPhF+gg178WeomHVsPqBxCoa3Mo3R1tpbvLSsC8O3TDiB0HYDXm6ozK63H
kPzKTHZsTh78tHICHT/Tto9BoZexfgyCdKjcUVnJlYBhzQpZnsp8Zw0co4kJ0qmgS/LoBPVcqSkk
9HEeQffquGxhFL+B1NYpyH1ff073ZxdEBJae26OZa6vKjN5C2bxTH3iHoN5teLO87FOhG5QGCPz9
LvG+hhA8b4WpTe7uwQrS84vM+r/kKqkQ3BlrSalHcU5XCDGIY0mAF6NhAdxlXL91/uWcjVxcXNRv
XXNlpJwaxuwTqkarPFVtTfaM6299El1nyRCHu4YLPZ6UpyIRfq4yByfaBIXkN3iOWMFAT3oOwgYx
g2yY5f4IqEJeRzXLkxG0EZp/XSd3o6q/bRpJYI/8wMVPFEpGLCtXnfdyjIurp669RhF3eGwaAKnT
ENQfwITTMUk59RrLh6kb0agWQQs1laxa+HL9qWU7pd2wNPKnBJhYhdRq0mqUkyPUHgfFbxY3ejUj
u7fM+KHL7LkcX12N2ey7BujGO4UzPh222lJF+dODvKgmjeIzQkd+QzGKWwrr74JxsR+wXwXRU+yC
ZcdmRw7rcafnaM4UCOlB/i6SVYU9WJcyyf8kLW0LlYKv/jdmnC1X9/eZsRKJLaH5ojion3q/CBYo
1lEV1KFylriXU3IEMZ9ibwBTQpa/vIVKti/4MkEUaCLrb98wmKphtoph+KStw84frcdn7sD9KHa/
486QCcU3qkKIA+lI4e9Mw9+bQRSSCsHkAxbXOJD6JYiUa3ROIfuT/bF/ECD/allUQCdTvKTrt6RN
Mhfhv24YKrgOfC1lJGASiRT6NhcT8IaRGembgmA2iKSTVL9yqweqoQn9uttdW1xgAeUCHTJ2QoyX
nx9rXVDJbQFIToydII9jBfYNRClniE/PDrftBvd5MUkE+ggAMJhlEX4E7oHD2CzKQUcFJ/km+dw0
IDNxEA6wHFspb/nJiG2KbPTil9V+CgL5SS2gWZjuRCY96rNllwr3zVFhCSlt81y4L4gTMrUCr6fS
1zy9ecbtN6Y22GTYykfW6Z8vWOoLk4tCtfWodwKmPsxi/l0RfDlttYNQqqMKvuse3h9acWBsiWfO
hJlQ1tkyKKGZ7n++DFOyqtzUt8Rq2fPVD2cye3lSCs0IwhvTgmsNDoouts6ZkrTJRzdQpVLvf9se
izmiqw2HDBNhObXJEqKz29KI9zojQ3FKdv9E/I7nVnPvZX6ry1EvJhqbKdg0nZSYQWdGeAbQXLhW
hEu5Si1GxXfKGyuhZqOoWUtIj2Q9pevTQAT3NXqiScl9Ko0Fa4O08ieJ/3Sfh3NIFFnp8VdkEjJs
BlX+d8kih8/gFrdWPNiC0Xq6BUWHLs7hs3XocMgIUTLfPg1e2sP8+JqXR8XIfV544aF4QamAykGj
zF6251Qcx3K7+vcZ3x0f2o4L2Cy2uaLZmgdBoo2gUip/k9ilvxcHV3MztTLshLstqRqXB5OkFRnf
dEe7UvXgQJaFStRTH6bCdKTVIUEmhfuWTF1B+kPFIVoC+NqkD6dG+QHEZaTWKEcFESVQHLPvNkkv
Qqa8foJhzqz6X963oNajsve/YdIO0iwtBVgBAGAP3q1lF79nf8RmufDfSJwJTu1gdPMJAHzlt6jj
5geKR8S7vyRvnPwN5VIUwWBFkQshVjhYBckf2z6CibZNNpLs+VtavZ8Ww+TBYgmz9xsIrJhiON70
XDlWJYMOY2YBRQppZ0cXaTdq9lvgEUsgNiuws5LjsnJtGkBSNQLtjnvmNl/7LONQklG+y3fBVK/8
4AnV/EBdVBdXPFhCOSoSjsL4W6qa4IvTM7SgBGHzlLLS3jF4AAGI/QiThkCiTy0FU611fl4Mn5q8
IPCIwtDzHSC+mFzHhxZwsX0li/3xn/81iGBgYP4fp1X+IEsuhpbuacPBC7fnxNbew4VmQHJ8k+Wv
x6U6OPtI+rHq7bBLVR+Rrj8f2mdmh82K7HQ23SGS5UQuFlejX3HaI5fN9zfnqP5qb0lXeaZSsl4V
+UC4j6/d0q5ua+uFaATRBIQhT3I+BGgekF2d3/dfo65d0s9+9FWZ1mXH7nG2yG49Oj9YoWGP1Z44
S4DsJgc02v9jxZZWtHTDdPFNFM0A/FnZ4GrlkGHykUDW4wz7ueRH3TVxFgD7WB1TNYcc+Mw+4DC6
3B6+MunFmxr+fUm5vcV2DzVjHG7zDiXErDwCqOkFKaonEztCetBrfSWaVyw8PYAYQspGHg3CTeFB
na03pCqIF+UKFQdAMvvDhbaqoIM5+/mPGEvnC2H3hWVTnRn5xRHSlV5I6pK1FdRX5qmFlZni5jyu
IWNHEmwxoubzY5z1QMSQgRT/F+nxZpCTFs8bDSsJqmQlupfX2oy3XseKEOkORztBC3Si3SaHOVZY
ZIdvMvhETFNwG6VDaHmwkUlX6hqdkYeKEpoWoh3GqgFYwITpr9Yex4ESrNVZ0GxxsTmlYjbIuqBu
L1cKdb7hTQqiLNIMAMsbx2/oHnfymNC2k5MHh8IlpUIPvvxeBVGmuwjimETePn5h2rrECXWYAeGB
NzT8ApJG8EBb5H/CW801k3G98OhmaggYcBdIHPtbeNwrjDvX+n1sRoTOkMztmLrRsiMMMLzL77or
jctEE2MwXT/lq05LDf8kdFDz23srRdQxSmCAa9odGocwtgKw4WJsC0YI+G9ZQ0NAt0hnwcMhZZ0N
YNAvDYN0Xi0ze5fFc9fd9Ymz/PEVsRHtOMtRY3yAYKYzAj9nbvv6prnEOFYj1uHKZAWOhQdl8ogb
H7FxmrDnxmUWH7+ZX79XfzETF9R37QFHDSIPh1ZhOHBs32Gg1xB8g+UQNl8fyOk0bGWuki6Njm46
mzJSvrsNL2zRTRjpIJCw8vcs3UvSgGqXsMkhOcg4IQ8SpEq2fSozKUMriCyGlNved1oMgxVZskFG
l98WgM2SvV0wtGHNQ0HNYea/CwEGXN8pRfVgcLeL/MVP0lD+DTuKbS2Yl5JpI80ul0rRJxmf6eZv
Uq4ydrmZ66+X6PKzl4QHsAYoyWxkkoovrcJduIOLY4xSzX1Jgroy98VOVn/0vPrBoxsH7aHsOz6k
aP/VO44EM0KG2d/ISYkITCNjcvUZpq7XQS9OdX7EetlUkmvFFiThA5tKVFik+BTdDZhJVhFA0Rt3
Eu788r0WYBnpVuSyLOtbHdjJfmUpZ7haKN8OdUJoDuXqS+5ZC0MNLGvYd3l9Fnm0Q9/ntpdVBBFT
zaurNyj28ILkEwTMrplQN42SZW3MklJCyJC4qXHm0LsRYBHeg/5H5+p6jGaPp9N3boW3WjjxjhSn
b3FreVwb/jKNCSO3tcawi63h6rfcGYFVuisBwDfxpFN+SJBKAUMoqJ3VeO37VaRJEM9DGq5G89R1
avRladIndhuvkbjJJ3ZTIBbOEEYG0SS9qTgpJSoTRNBZ8SrQEps4zFunW2xTDaB7nM+hMsK8dQHH
63RBFzDJ1RrwDvLw44pLEdl9uddsqYZavgh0BVaYoPsIIYBihvjrIkPjRM1c4M+ub1ffVIzRROTb
ispC7G7KIjTsFYKvATM3ychFXKmLkK1+67H6+7FYN1VEybSl5lfDaDkmZz4QJwQgLo8aO2jtfjDM
jray2sQpMomwr7cKE06xW1aSnND50aaYyjjwk62aLoIavx7EdV97ZGe9fKbc1Eb5ud5GU7ZSVDEt
guxWuq4M3r8Bq7QnyIaJbxclcuRL/8ztr45yampFcoFH22Hvr8OQqrUnqTH7YsK0ludGvLxMtt32
7FE9qlMMq0F+z+pQVXNPt0BSWy1ebmmNv8I8xwVAv9nTf2Hik3lOvIec4CZsJOioqv7DpRG8f157
nFPH00raPYJPkgYbKkJBQC7XEu60XoUXWWnGrxKuorIkjETjbkr8K1Apoca+5Y1yaLm04UBb1HLX
o+sCg+MmRJEQqGyVDYlOAQinDsNBBEb0njF910NJ9oKLknxyn16PeY4JJ+02RHqcVKq5M0uOOQf4
g2gSIMGR53zrCUYNxVcWsE5EP0KUraUOJxgQXPWQ4Gv/HpiWpiGfOsf2DFPK+psz9kh277zqZUps
+9/kEjGpuhIi8if5Et1CF0QfHFfWz7GHPPE3BN1ifQVLtHYyLlCrnEsSaxv370vtLlDths0KZBU3
igeJTUqUldMbQAZi3+EJYYiIlmj4VcVF0PC6rz92eKFr2aBIdwI8mm83xUcYnpHmzSHzBCskJOJf
YO6QEMkms/C+joZyWC+Q9rCywbiwQhjGEbWGr9mLbOZMlk91ov8dI2enzO/LSRiII91ucy5Ad6Nv
5yB1RKxv70Bu7xeqABlpGnPucWv8FL6nY7/9mTePUNljuQd9MTLrwaoHmtltKtNqhFS83QmXo5Wf
L0nf+Wf5NwKMHPh52lX/RDEKrQNKUXB4VjC0k8ADFgeRLPBlcc/L/YOUKUs6iARfjsv38TXREKpm
odnLv4vjvzP+XEXCpZ33fpLjIok9jKTjqmVngWzWBdOod5D8yGqnJaF5cvVzaBy6v96xxS0ooQnd
Si7kbx3lmDaFERgPWnpdiBMhu2p6e2uVwzIJLguznoVWLl/ekU3SW1TnMeVL+bqXpGPKbDZ5JGK2
dxcMoMs3jmgiaTfQiaN/YlwSkMcLV5O2X/uoFO0Xrh7HWnABsk+zbvHj7iuxjhXjGQc3ZlvJAGwV
ydVgYkrqU7R+Vup9aTPvm0dhAovyTThykFqQccqkONpRxvnFxsZVprV9W6FFwivN2vK2+L7WySFx
yq+PqIPLZRvHJphAQp/3n5xhsfESs9DNrJ9pYdW5kiTQzoG2/x/LGdUenjsndy4z821F9ju3IrWK
9g3pu6iNC0nhFN1i2Rb0e19nwsuEPGNyQmiACOyPduMJPKKPFCqDEdw0IQhXowpAk4OZ8+DjX239
qtG/rxpJfA268U2MDFeoW70Bpzxak9o9XXYZQ9HswZq7v+gZIV+gxiTeyzFG05ZyAvX5kIc4frP9
7Po1017l6wiEukQdZv4S1VUwiHQASbmeGvePIh5q1q6z/YnPLMPl5txWW7ydVf7ASEna4ESjlCG4
irqPkazAoQGD3EXJenlunmkQtfVOOoqVgRSzEeyfbrskoc6EY9eDZ/wlM7T5luI2xs4govIT0bFj
L3fTyrILX1ZhGTjDn+jQxhU12ZqXhcTEE9sCgMsg9zGUB0KA1kr0BXghimhm51PBDgGgyRoavYTF
IQp+zkLIMGSxsOp5Klk133DAgCEwi56Ztr/VZOgku5v58IifMVopWUc4Y3owO+rV+jhRgHn2KItK
axtKcDLxeWRXpTyPFnIXhJFPP0KT4v4AtrBvgpmTjlLtlnse93al6tjPrdRMOGiWd/ekEvDn1MrX
dIc/g7Ao3yNuUyKrDFvwJYxJCPmkQlqgElrYDpkXt3s1AkLd7HrFKS2R9P0q4EPeDn7MS8DiYk2f
Aj/A4SXu5O7OOgWYu3X9yamPb74tuN8cjKtIH+ve9r/GUVOYMmlAsW6JoMePY2iKjV1SKrJcUS8f
EE6ruFA/KftXXH4hViJbL5ZKoFhWPc3kMjYwkjLwgQPhlCHcUVMka6rE3KSzo1m96rykTnlceHFO
GfNl4xmLDNdru3+qpVH0KxeO6Ib3SiQhUg4/gTfLabc1F32+Y6PQSHLn10LHAMDtkktqZ1QS1Yil
JpDvXubIpvHEfQzHM5dDeGzXMTBu14x5+q8s/1DU2C+Q0wott3xiIdchpuUH8KFaJCGdNCPw5Jo/
pVoTpBc5KidYMjWoqCMRs0NGxx0o6+EIP0z18Ng1cKIumgTzrBtQSvuXs+qAEFyfCtzxXwDlg1b7
fM6FFvwz88TLvB6d8VFKgyHFG5qH4IoKdV1Sd19GmYkYbCff+UjKnBa4jJQ00wjJ4VXrPSgngLYa
9itkpz7wBpGJ7+lbzEVWYA2AawZSsKCL/ky04IR2qnf9YkNbzT3F4S2MwoJNeFQGIOI8awcB9mbq
p3maEV3jSqEMO0PiqkwfsoNyIfkSRmDxD/kb7Z//5I/ZFIPKKclVaU22dUJAIYmsCOhOa1o0PGh0
32xlMirvNlHShkAcoyx9NSY9wRnfK8pcpAp0edvlU80q18yW4DIA1UZYwxdn6ftIcsKAJc5FFi0s
6wzRueCEcKJ+wdaGqMJX8QBqTkc/5q3vYjZyhcKO5cdFN6nmoQVJcAgJxIwkmGyLH7uoj++eJeJc
UBzDKonLhyM7DsRhTwgB09eZUwU/Npj8IIL5B1Hzaa7ycFEMQldmv6sH1KsKWzMkv0qUjciYpuPO
jTp82Rxjbs9FhHLSh4w9d9iQe5lr6GUG63qu1hhZFntAeMf76R/Jh1ON+UkOaykG7ivrnrZJfrRu
b1L3Uddq+z7B7n9mteEJ74IbUGSB6llG51iPGth8h86zdOq1kwITZfq3eNLa28aOEMJhG7DyW/gt
ptl6qeP3PX/W7ByZn3Idp0YXuHfFty4/KB0CAsWjcvCweXkURzidOlEzahkNehz3oUW7YheJo8Sa
7iZyMhZmx/XvJg72hoDT86u6TC3Zn02bOpbDjEdWZ3KUBQghqV2dFV9tY3asxwcyqOduyodoep3t
AfZed4ECrsqDS2RtV1DOJcm7zehCLX7XlmwMV7VWLVmbEEnQmHsv5kBXelQQqvGigIdOEUl1gKfK
YNnQ136kc0v67RP8zu+Q7CGHi5RXseSIN5V7dMI7At6AlSmpCfw8kvjYTVDscYKD4eeYC1p4MNNM
BVumgPu/801TtZGhOWAACnAN02DD2PQx6HFy9D05DEGaa18K/ngz3jXMDo7ci58NbsmxMpg0MIio
ULGmkQ+ZNIIayO2XtfRx1XFjHB8+88H8th7WEKhpueUzG0s9nairgEjzfCzA6PopYebHH2XEh6UY
FSjP7LIakq2tEVlRkDrApPvT2DHVJeIEANJ7z/takFKNycqHwNuXwkl//QnXUyLgQn6U44ILYK4Q
Vie/qoDoysPscFW9titvVd56wMbegA2lmG1rg3FN7CgMbngYrE07aS8CwLulpOZM5G5zM8aApzMv
Oe3RPuYLAjzPMzTdYT+BGsvGOir608nUMsd74iHQ18w13W/wTx8ufh1oXdP6U75cQ6MODkZwrIXi
CchNLYYtE4vt1J+KUzLFf8oCPN1Kw6OIjJyb3N9Bx7SmADhG8SEGTesJSIM+NZYgxMKmatt+Sbjq
wrf/WnLTr39VBLkdV6L9EYEYwGVa4Af+Pg8V3iWQlkE+6KWczRMoucMJxbfPBPAbhfAhFs/EOIWd
jtpTBhpXWBiRH+ltnVyoMB/kV7ieVNN8ESTbds123UvKBUSfv7yU5MBzw96vv6FHB9SFKRKC4eCy
Mo7/qsl4OwvRYQuXd7+zMPLbKPp3vOvEPB9vE+4ca9eNSo0HQpjE0sYqziicxrde24G+Nf+/S7w+
W6Mcv4l18oQnLcln9fNCwOqjXPJUoAUq4SfqzgdxfzXCQL2kbN/FA/0IeD4UCohK2ZSzAH1wBESk
SwVpo4n3/+RSkrqqcnXYmT4PAgU937HzGjpUoA5pkRsOrv2ST+xzia4eUpKCGRKAqQcbcTfBOZ5/
FmOhS2+qVBSmKFEzmkfIJtXor0IxjcRv0CxKWi5Qqe0fMKhUkYDuB8tqzYGEz63HCQxkcbHUBiOZ
TWCVdV3DLBmXktslayKpZHFJQtH2xCYrecAouyg7g61qpMq02Ug1jM7AeOgylCUx/8nRuSHm5j/B
+6+h6jwRg/rY0R4iL7oZZZX062KwDOiqORv3enxQaAp5LyOoEySHv0r/m5xxXYZu4a64FRmcDmAO
6veLbvGFd0HJ38CiDiW6AmEnKD4Cr+EvB0ESDWPCWcHURSpjHzWnEBOKXvBE061m5VZzmmgjEsgi
ZlW9Qztx0zzkf3LUpXrKYKhEFBzBUHCOTI5IteL74dE8sLHbRvKyjPDZDoqOKRzM9GLJ06Bxf92z
VRN7IT8v4bH5WCawyMEYEeW5zsRrWbK6JGy+Sx2mPIYJcFkXO/AU7e6ZrUOM555Wn8yY6L9gZiD0
KvKLTtoNmJU84TZ1lV82ajrKVdshTsD1foDRVTtUWEM5zikLsKnwIB1biUYr68YOH0s/gSjDY8JP
v1EuNs2OR/I16+D8/Iw6QBgqkrCOSE5+RCG3BKKQ0fRU8whI3sIUJ7f4INwXT1TYgVbUKYpNX3lC
qAZLrF5ooKpvgLm2iVNJ/aAAf8MOfQTVdmfJ5jGLKfgMmLPcuzBpTumndleDB31BuCLUWv+1qfp5
LZ2rdGM0/2lDn9zNb/JDKtkUXkcZY1Mpeiq8jWbqfI0IPdUe6kt8lYsLDIua0g2FZ/AYyDFt1hlM
rkTMOMX+ArR+lMFaBi+1IcEezhcFuC/DEuRG8uzSiHe4VC3OpX+k6GCTiUCK9vl+yaQof5TtMmro
YciFgdgS5SuTQ4jb8YB7Kjo8pPntcJJEP5NCT40kOlI3RnWV6WOz2DCYhSyUDwB3bkxS6OTMAX4t
n14O/DGTturwA9I2BKXrYBFx9b2xbUSp9GYeckC3avZ3aBvilqDwjYFNJZQFKscKH2hTw6UyNN+/
WIytTpqG3lC0hK6QH5QNcBpIu31nBTikcekKBLK2skzGD76ozD6VIRd4UVHX4YxYTNe6FuJz2POf
MUF0m9pO0faU1NRJY8ZE9Fs3ZSKvS9lh1D0qzcZtfaTw8kuFtD9zndlcF29x9OMKhzI98oQExilT
eJztuOfOHAANdrKmp4ZVhJqzsbepX416vvWTHJ2Tn43OxBXBWkAfk+tsnILq6KVs064cJbOHTjrs
twjqNJXxuDPMHw/Ef7C7zVVfHMx/EAUtHQ3rO5mGzj+BWjAIZpaDVzfDX9wE/f5cCrRLMNKDpdg5
DlbDedT1D0SEPNfw7o2/sYZW4zAk75A3CmheKE/AG7j/yZp06uJRrngio0rMdVsRMcA3pauObUxw
+0UX+EEFtrDi8kkjvnGWc/AwNyXmeLJpvqPgkoheWLUilAOz8T3sDFuv2dezFHCdA2gY8N9Eya8m
OXeyvNVKqGiQqqbU/tMpqwCs6NOy4xLTz2ErcaTR/cozUBiyGZ4kIr/xle/TMThMobLjzMG6jSKv
Y3fNhBaeuUQqX3ufXO4IFMU1+zqTEdCcORMO65jHuymDZctIOdvLq9XxTqR8pGhAPGMEXRBl4BL2
yst2C5N3+aiB0yf98F3EJEUhLHtionrdd7p1wBpaNII3drB2AmNQxcdkR0jJarSZwhwOZP9W/qGO
TmXy+nKSsqWWRdS+egvIkn2HAcjz2Mx9do2wKKCMxDk8UJcciLsuqaJpoMPz9y+Quk3sPC+uY9Q6
m8gAbgIdQM9+0DwYWgrx4rEuxdOrR9iHqYkN1Z1ASKaMUwnzLuw+X5bmCCmggabovDIwp1B/Yo6i
KKqDYCTwdyNXMl8V0vqKd8lj8jjAaTFetZ0n3BWyH3aiPYH7GKKm0YI2NlW/tqHLW7H2WaWaa0Iz
T3nyPGE7ExbH+j0Q9otLPsd7eXyVbSmcChjntlfguhGf/BG91PNC6C57MLCOWgCcxvbfnP7btY64
kz39GsmZqS73t+qqkml78qL3nqiNpRy41Yccq4XzA/8ovhhzGXIab3slV5nB5Gvg+cFh+HHqcnAE
V9BbwgWLlWWSurbZFC5WrvYF09IfUNTHU1fvkfnS1wU8yeEotraVMk6tgET7bvoaUE/O3Br+tRAe
BccQlQxPsC4xeNP9LMSqH+k3um2E/Fd1UWfupSfKwiJyWcxBCpMp/XIrazVgSgefhpe0updHFWOJ
u8VCScKdHsdzYV5bbd+8zH/V84Pr+RvWnmFKGJyaHNKiLXvfF8Q/EihVbQ37//k/zgLNpmK7rbUm
7FGKJD/ZzF7Q/oaRvnjeB/LDbDoEA01nDYMrqeyM/8ZIuFzNmoSz6eULZq0ee5+/f9axfJAwuTvJ
ZfSjaj0aPkxPKRUzfx6zbhwuLGWiLEowFnDkwGw4rtuC9DDbuEKaeGOPtbkSNbEEczrRT07YV6KM
FNoYLNgi9vbtlqm+qbulcZ7kae4FFrUsB8FJ06zRN7zzIsd51mIUkYvMMpE6TGOrz7kLuZ59yu5U
Ts1XU/6WOH8C9DK21EuWsRPOLOG5AyO3IJR/nwMbjQeiM1bLDK4UyMk2pjO6Rkh4KsKD9Xz9MFG5
zJx2WLERI2Fd/wLVbjVfLf5foHm9ooZP1v04WiG/yZugqmT4gZiQPLs4cTVW2pbKMLlH622JkPJC
1MutUnhE/ytYU7/ViXQkHLA30LUB/J7S8N7/KIBmEUmsgX7JtnoR781tV/kYoxqog8/pTNxX3VRX
gCHrDrZemd9IQNU7o3YVs3xlv1f0n5dUbCHkH+y972y0C/CBfZgDfSEcfJkh7ZSlSxhKwUMEJaBt
kFNLciDEx1BEWZMFy5MU9tEPCoowtkGVEkpxHWM7vqwwLduwJqW1WsPXQgn51iAapwPSjzxwP72n
BorKu3cvCPnb4qdeqUXe/XEzEyaKGJSuGJJUSRz/ZXgDGyVOA7oD3/DZXv0B8JeClbgVyaFP1sOl
c011Yq1Nrsn+ZzWe8H4hRNlBgGSu7xXlyxDVwbYbGYoGtll+mN6LKNemK/Hbzsf9dhB9saIUfs7e
9wzvvGzuK2x2aN/N9xuWWIIV1OPkynDmrrU6dISf3xwe+R/FM8UNvOMsCZ9Kv7EcsOV84ZM7eDAN
RtURdVGYMaCLwDG/r/41czsxu7X3U4YRQ8dxSKXdsk4zHkUjEIrZsu14KoDcFRgMgqprwgr1G1O9
mh9vQ6qSqSMW+vUrQRPfo9fy8896m8eWPi8k5HQlkn/TwsWnhl9NmHinXAPSuf3Rc21XL0qCOM2t
4V49RZmE4Y2wZbEXs4eVJ+wg/EjgdQZiO0XLoqcE0ddD0JrUvczIfWxc6GVq84LdoyGTppdMAeSj
lcr2Cymc+rnDvGSXLBx/9FyuwnJnW+K6PI7GKw0eGrfutZL/ptQXRzYPMSCucbpFecs7s/OsyVOA
xpieDGdHFX4m1rZIaY1uqjz8rzR0oR6cKqRReBfpPTELu8LabrY6Fv6Q6ICdCZHhdDzl96js5np4
M2QFHpRrQcVrUytBzMpo2Iwd3M0EcuoAuS1VJQV0ikoUkj7nSlr6g+aESnQj4/0jAiXe8o3dwh2j
Be8I4Ts5gTwrE9T9UTYuhquFaactgK/bUPYPfxij/dfx1SCV+RP6qcQ2Yufq+jFx2Y5drSCDYK6k
C/yuwmh4geEHFHy46iub7VMZjCdpNkm+5SZtpb48dIzJSmHj/elOZ7DZlB9sJCdbB1tnjoslP4iW
tAkvgfrjoDStqToyVjDPWOB7TIKeRaIbk6zcREx28bOZkiL2Nj4ZMfScSXh6ozmAVfTwnnxB+8xu
bDURi6T7CanQC9rri0aefgdg7RN5KB7VKdGc98HxBVz8HU2pnzm+/FCh9ZOmdcGmUE1NCZicLQ35
wuSY8i0GcfHaCOB0yeKdufq6NsvwogEuAeKlXN28bg2dz6RTCE5wnmPRQpCSq9GzIXGL5HWVsyQe
K4Zq3YTOnEdtg6HMo0IXYGzcK2eekCu+rGrTuU80wFvfKOlhf9FrakQnB885jzxAnc6ybGsmZPLa
NzJEGeHXRWDq8HZh2BjQ4NiKcDcFQbRa5kE4tQ7gj91PVhHxjQzhCWml9Mmyk894NfvPn4R6YuiV
1Gc8IlfgveQ1rqD6XuqGu7No7tfhBGvakfE0OFTZIhiHL5ujk0Nn8rsnrZcpzF08huyEQj1skHr1
HJS4UXLre80YkzQrpvjS9GW/tbA1S3/9m6ucOw5NrYbPhTKd6/0cb4dGI/8Sb/WtrD06a2aVdTyz
Vihd/qQGB/NDE4z2ZQ8y4Q6SeaWn0pLrJbZcSl8nTrKAWL5hokX3uDCF/aUPSzMU4mnERv17MimI
w02qlxEyZMYUNb6nfJAmKaYN8/ZbUEPQ+3YxXds6MfvRo51cSPChatfebcli1D49aal3HNxdJbOL
ySh1UMo/RhAkE9ddcAowTL/hDd9lIiTw8nrEQeycULpk/weJKiEcwveC7eSbjNKc2pHRe1mGgjUI
BKfndcSCEXfkOvorJVOUiQv0bvaX0g14K7odku6aqcnWwC3Mc6o3xtlxg8UrJXsvRSgxur7dJkHl
C73PdyE/tdzEqzIqSqjZO4v66vg0esNwyuuAUUxpz5BPuiPqfBXDjwhjylo2uuJKz08hAlvHWv25
MVNzEiHQyC0kDm9WNQ4EmzxoH2g5WM5U4/nO7b4DfNv6VYBIeprhx9alQNYI6z1IYpvYsa+E/N8A
yd/iwjWBlswGhf6w0noV31SkLPdQzOm9tPK6/bi0lHpkq7q7p2Sn+qzkiGN4g1z9umjkJlJ8ABSo
rH56TpAERbucKxnCt9pPUpDl+QsUbkefS4lZRCUSHIJJ0mcOE4mFTlJ1ndTBCumGrengyNiwz0PV
ynmVfhTHgZUplUVfbhxNaSV2DdelsSnMOrTd0TbLBwehWE3Nup85zmfkl4UBCN+68ttbuKGVVc/x
bW2Dr7USv4vOq/X5mA9qsCmYy5XbcEnl9ugmY/7wuEHArfMjoaFchcgICorWhDYI/VFPuu4DlsTX
sQLcxcJOJYHkPhXRivejOA9nj4U54U3evEphxKUKnyzMY90YO4ST0zdC9qDa7f8ZsRhLbv/gkEvp
abTGSA4KqiWy7E0NKzS4j3lmjJgFCDingl4X0XJsE4HikqAEkjNWlnp2uLzVtk0EXraijJ54ldx3
AFvW+XepJnzAgCVXSgq/qksLAOFtAQBZkpbAblKG8A4e0ehUScH3ttFq4Ojt4A4htuWD+DLeUcAE
D9Rj0tcpUhbkaxIwaHDAwC0RDpMyhbiINpVPmW96txWEYdg1HiE2f556lAzDUrDKMfuo/eHy2BCx
q31l9IXE+6+ilYk1SFCdiGCzfugYDZlQbUtDhe4PUsGi3hkB5SrKya+H0xZX1zMkDZFz3btYSpCf
Pb07yMq18c3pE4lc0y2Nckb1FFuZd4tm3zCr25z2K6l3pFDDMH4DntzNuy1gcjDoQWFfqLrL/gqa
i27VkK9F5lbyMm0HW6nL/+oPLEpsF0zYdFu+8PSXKaL1StWmn9noTTyVyinkoopMA/SoQAPo8ZBA
GVRibxLfrr2eXS9bhnw5ymzxBlEAmBS/Cpl8abzvrH2k+7TTyp7gHGhlfCoRVsK9KGS6j0BfJ1ia
xVm0478Iovf065dc3pIrHe6XYAvzvJhA7zyTyfCHtF0NZJgo1jaGf0EkaDE9PfiSF8FZe21q/QKl
7Qa08jIU4PYYvIAs3MubauGyMTjpPM1rMkgItWph/nyuoMJtN9MUAnspIYlqfnfGT//P8/0nz2ZI
vn1vRiLNwA5dam7ymQxbn9uqGZzVA0v0HUKvjpNOkIKSdwzfdGWWYH9ND6/t3mYUB/tJNZCLp9M/
Qe97S0xBqPv/WoO8fgBLW9wb5XUPY3OSwSo8cchUExmCwLJmr4UqMz86/paQhWEKfvpZbX8C67nD
OL6kyI5LWSKK2TK5X1H0Js0N7PQle9mYnHkVU1ywYaJ71n11FGIiUvdsGH6bCDSFOTNlnBCfDdUF
CExnPQA2614WnUZBf9EguluL/jKk7vXxLnFtw1kRzmmW0UfZYqe2iaKk42GdQXx0c13ul1lSf5h9
u1qxcjDSKuibszT8bIHthcL9/LOdE1kfwKNIS6ajL/lngzKOabNq/08LUcGnWK0aGxtG/IcD1p8f
WYO6OwR7nBMYKgUpl8+Uq/QVaWZl7FXdjYT4pYnZiP8CiTGrdQOvca+X7rXj4uhlw85zXcBYa1cn
vwYzdZ9Ws9uEE/L/Nn1mwCyIFRHXD3I4e9k0ADOPTgEq3kbHIZey9YIMKY60k1UF8BBCQJZ7pBT8
xjcZmnL6oVQNhKwne4uYC68CEEgBKgkyQFliq2k5Mf6ernweL76PsdABLFsXUKDradRQrreGenZs
cLF8ARp8uVKh60Ai0L68NSqF90Y+4l2gplUjF5UjMfD41sR5N40YuuzCuLDIJBrO/d0Gg+n67NSa
3mdVXdmvtcq/hWwpbXjdzhcB/r2CYQoY538w0Vzxzee7bhMeYVBJdeZgpmZNVJi6QQfdAgyrghs3
vDATnZDh8zdBWUl4aW2SAb3ATp2yfngumlggNxqhxXI46VdY+OsZGtFdTh98V3/enKY6k8DpFDvX
o8kq4/OVMtIeU3H14Ls0zlQyn18pQJlMFYTW5/bJN34AUhiTOGnmkOuxYpKFD6clBP5lY7w2u1Fv
WFaDf1r1xL3qvtzVhbbVOckDD25FHqtIO5HC3hKBkwPiOObIPvmcK46Ede+sCyaSSDcIiP6bFxdT
FWK974DXCCQBFwm6X8s2ITSUfrB3s6dABq37wuuCqED8JImYc19+4JzwILQe6IP5UvLTuqNyOmPG
cOorZyooRHYxc5v5MoV/K6LgxQuk9XhlICaxGcKApBX23iy7G4VGdqMQp+WMODBvDsplwjOakc3W
01a8sfYyP9w/YN//iH39OZstxur8pfnIKPWG8pSk7XAzsNgmO5hAoBpOPgwdZcK6xa5610JqDOiE
BxtdcGU2CwfeobdtkKWNPtlnWt1fS/k21Zk3feg4NhY6OzjjRWxT5w+0ZlsuQw0XnDS4m/0T66rw
0lrHniBw4xMC9NJFDypEamPAojptEz14jUqbCm9hKeWh5TGWMk9/Rl6vwhi6mrxsI6ib+VYVvgAc
IyccfAJc6DZF06yQ1kuUthCGJthaCC6c6ksspzuIkCzno26BdhTruOiK6TJSg1YSpi+nZm49dLCV
4LVI+xOmauy2Z+N4uNOLBysTDmkzrrsZ4l97+0q1PzSMYC3t0F/3VIwS6ZsTbTJqt0Q+aE736DtL
/nw4up25cj7cVs27N4eGlzTO0gMSFYZsW0/380QQynxCu0OpajhCOT6PARXYH2KQp9sy/6Z6oa8G
IG1yjCqwSWqq4g4saqNzgdpZveliPbEgkkoW0nxK85gfavczQi0nCI+7Ph+9UbOuQ/879Ex59Eml
9aYzRFUKH9iXgPsHbjqhXfT8VC2DY/KZC29IyPR1c5ddW2Q//2bzPOHmYTpINjtgHLBTxMxhqRtp
eVJeZLFlLqKTkjcbNrlTTVy/wLp/f0APxpR/d1vvD/LHjjdVTPlIAVIm7SOFCqwfwKsQQk+OU/s5
fabS+hdHD93YtfgLNuJ4ieV80qO6H04nGmdsLqTr5ERDBW1NmRey7e0JMJU7XJPl5o+ch9V7a0/K
Kolxs4899qdCWeyhmgmNPdMEcpvAq2vybpW9xNrjQnqprKZYQx8ToG9Up5eAJCvFIfWWRKe0kXTx
FykJVNbmjeYyR5R88p43JZEg/nDGHWJdCOd6TEs/qW7dkED3Kwa2/6FPUt9B1hb3Q7C6/VJ42f4n
rxv30k0l/26WQ+VZQ4dykbnvi5nN4tt80NLVj9S/g42Z2NS3M+pftQslbNkh6KkQGxvPE9JLmpnz
IoTzx2N7vfZ7/X7DI+tyHWXNOwA0oMr4YCYLHVvWwGaxOfgQ9zu3DIg+oIMKRAyVhBCnfltzIBJw
+BFHbKWuRaH4C4SmtijHAyC8P+xYcrJILAEcwmPPRCLbdueMt738mtddj5IrpEx+XgvijoUqNdad
EvK570yehDMo1TTt5QInzQt/p+eU2oJKYjlO95zrsWEu/ygVh4ufwHpa6i3eZI2JjvhEInJtmf4L
/rKaZRdjVPybOrl2UN8F2uDwKg2ExwW9TI1aEkCJTfVCIbiOt4A5Hb3FGu0aXIRtdfA/ZZGFmEsZ
AmC9PEPoCQRAPmG8ldZncG9gqC2PFwOcdVF6rj/p3MNTv05rznMBU/KcDO/mVeUEsh9Lf8kQfFCi
phfxEvenZ51EjJxhk4NE1aYcEcyLHQ96PftfnhALlgwmaOFQ8ciV0kO2QoakO+LYC8Zn1oho2CBu
J3ZUXE2HnUJPgeQnxnWXdB3wTpG2nf4aU1n1KgOLNxB0BPTIig44QF5HuCuQ5lv0/FE1I8BFkQDo
KDiwCoGRq2huwEVkNxAmMsf+at85jBLR05pg0C/i5KWTO2UH7Xo0QS99J5JydPSbhCgkcwQcpXa6
Lq5U/rPbzwIhLJzX2P9pb8HxHbX491amwTnAB+qr1fIABidNsjmpERS9GkWEtAyAsBYdWzUn3GYj
MDcxcLtgXrL/zrqq1b6PQFkGeyp6Qb/D5ntSY3THG9AiW6lQRoUmjRY77g7zZZQzDWtnvKez0oK0
DxOwWY0inJLsejyVMC4aSrFahw7puASwstRYFzk6ls7wO1N3Xoor89MWSQmM+rWxT/tYDmxbIK1Y
zY6qRw5R1K695ef4j50N1uFeOyY/5Ul733Rx1Qg5Es9Wlpf/othRChC4OaVqWgu+cfnTwWbCgQRq
ALoB9czdGNDLsEd+0oJH7MKgeDCygNKGFmFr0opvTA7/wse0xPomG30X0CezA2eLGogUyBtai6UV
Ub66lgiGBe/imy9HTMDKZlQKlY5MuQI0wiyuVzF1X9R+Ro4xR+ibC9hSRWCF7XdPywl2OEegiqQM
ZMbN+0xHuBjCQ8DsgVMnf5rYz88BKPUyg76IhZ1bL9fAgd+4EL5vnP676KyYF+j2R+E1Xeuc7CPd
fB4cEPUaArftVp0CUupELlzseL0BvQskXNHaYAV/fj0+p8bfni7F1D01kEgBR9YLGlXNLsmL3+IP
NvDP3JoQKzsKxKqRnD7qsOE2zZeE6hEXmiXil9lhGuHxsYoCoRK0OW3g6Wk5Bma+VdvqUN3eR7j6
2COsUihpFq+/wVqLfYZUaU0HMZbnGYyfJQrLf8+xOdIWtA0zUI/Dg3F1AOpnbTpdNIX2w2XNBUId
RJOGlrrQ8M0ndyCeAdarRVtDBWa7GYf4OC0lT8ckxd2wIpfdKTbetCnZAOUqG6651E060GCw2fph
DAPUREeABdhbaW8rOIOZ1N0jpiZDU/PFkM3pOOr1+MFLTgF7/05Z6K7B5shtRT2cCZNd7HGCdpsS
9P3KvcVIjG0c5L8wpPt11EmLwc40cTM6HM6PjVn/vh1mIME++cNjrtuZAmwI5vC6Kkcwy5k0Sm9+
2XHPqLaEqWXx2IPj/zJiIVE57gi48RpaLS3abXh6o7KfyGfQ7JEEN6iGHlrslq97nEnWUNtDnqAL
o81YHNxE5gtHsw85k1KsSQXz/FYRgvZNSrpdzcK5vr7sxiUGoMgn7O74Edf/JadvdBX1e+k3JSE0
ofvab+YTQNzQf5KroFivOJTTcuBlBK/cm4mTCI56pmiarWYKE4bL/ITrwPlM9Tjs1U/hLF20Ucdq
nGSfuxG8mtI5Ay29k/PJnd5Drajm0JlVzFmiZbG3DpjJ1C6YTedJOorRtOCqU1DEXjW/HxYE3MYa
wcNgpTTnShI0R+LZoG3oXUvhHpUGM7uF2W9Bf1n4n9WX/rLJ0wzyzGCq8+8DSx4DvA5cURrcPLto
qTYAtakVJ/ijx9PPMtWs9RAUGQ2eIF2K1MCe8ZmZozIyvhH8CHioFdgH8Kl/qsI9bFpRwvSwCd9L
vg434bDCqnF0o+KiISnIkBi+UcnniYKjijDiDiY3CfCv+/+wykFDeMOJAUM6natdP6KiC24IQ2ld
xd3nFyv6OG31STHpHNhtP9qW/S5WqwSwGNA8cXeTgxLdhRWIRKcax3SfBwzMNIEJeKkungB9ogkw
73YiK6qTc5Wi4rhwloa0tcSxx7SAIJhPvZl/jBl8CbSJBXE+G281KMnCxelhmRTH0OlZzBFT7xBx
YaOACsPAd8uq0dSnAb+izGQJUSlf5mBJNdR0pLpebLEeYBb6zFaZK7VKtD4PrvIu16UNPbzOhIkO
E8xfzwrkr8xZu2y7R0hZgqeFFR12JWpek49uSEZccAvJsLd4APYo9Dhon71z6NX8kA6NmtPLTbT9
8Nhvg3dPYhWHjyGbhEOw6DDB5Q84eHjF74MoygfluJZCCo5Pao6c6DQmMqWxbUs9u65/Csjtvkcn
tWrRUCGHIMfFJtMlI+GeRsNpGiR29JOnsPGAFe8YZ8qFrG7ShotNaqudbhd/bPGvbF4LYX2CIpv8
UDwBP96i47I5c+hRx1vDno8ybOSQFw056kUlNGVtvY9MmVuQP4/GK1Uq9NB9CYFid5Dp9BS5KZ7w
ZGDvet+gfgjSK8f7Ex1HAgE5mdWzMK0arkyE0nz3+Oejx3xVOZPyp4CXn2GCqvJBxbiz0dkwc1yv
uwteuPpVnV95h5uHJskPvo+o+E1IliCttGxXjLdcgHaehczEImdmg1UJc604Pxew7ik938MQJImr
tdMMHpxPaJWkXBAORTaNl7LqjEdP/qqs6ptTWDb2cvxlQ7qOh5S+Q4dXRPB78nAITLEptvU7VJoR
LzrByF53AMAcli5OFU/8p1LqFCSR4DI2rJYG9zqd+XPs0s9p0pRNpz7L5t0snQEWimHnP9TblNns
zdsGj3lBAoslMBCGBjaXx1uweygrDGJiNDAX5KPSfIGMD4h1RKkfrXi1cjHBKgCR11qpP3EiGVCb
uNsaNob8xdUHmdeqYoHsHwQmCJ9HW/KpdERDpcX/dBMo2MQdo7LKYhYCW90VPPL4Rz4rYx7FQIB4
QNWFmXWdceOrN1UAK+Ntj7hpBZysEJXEaMYs6l85hBi0OMzjWpy7opXviyxyWfz+zDovQKaINeW1
SVLrfFEylK/ddm91jrka7W3qXFes7FcxoBSaGxisTupeuQcKFC1I/Bqq4o6FyUqbIWubeLqfojrC
KNPP4duTtUyU3Bdc/kUK77GQozLd6dOFWi1PTEhiMZZ1EEmncwzYbBac+863oYd7v+qHCT38bgb7
pZjwxt43fYyo3j1fwWlZR8Ef0VC0ejolcJEckMSjYxMoIhecYktrM43XMgTMYYNy0udsjhyRonRP
vE02t9KZ8XUt3rtoc163izyj3Biy3BIx7vbTwP8p1G0wsriaUSnFwKHfPnbeiyfXANZcYcUcTqP6
B9xDJDIum4k941XMReoojSXNBrn0Jv6BqokTIcVQzfd6kwpZTj3aATk6Mw+W0mSJ5iyrG4V9UDaM
dJCMGKog56u0yG7Q+U8CMjrd/pYpvGM+ODpzDgSLEo9mcolJ+EQnXzKu2CZ/c7q18EmakLeDpAVf
KZmbIHDlj6h4n1E99wCXgRWPkwskFsPNzc2jz0xOeqXP7dP1/ymIUYup2Eqra+ra4QCe2YrDQ+HL
vu2JbAiKHo0hu2sXCgzzpLVuBXsY8kPAOQtZEAlqgxknOoRaM4yK0fFXRfkmluScOODQuY588Go6
77Jb7/jWxUgitG8KVm9GSqzbNIN/yzd+OYXq1BucwXzdi+s+gx5XoBOkPSEyP7uRv52itA0zWFgD
EF3gJh9b8XOdhoVc5TPKzTNvmDTEKO8s6iJ7aqho5lfMagITzfxFP87PwTaGY8Ppa37t6c/DRJik
/zq+rsQlHVLwKPuHa1Qz5hSVockF1fqma7folPcTLAC9z73Y8BuwtzikVFWZr1ZuWa1ycrwQ2TUT
f8cOQPvANrRRXgM21J+ZKeSZ1G6nQiLlMPVgipSB2U7Gn7jk6KwScGApLHbomAbkWsOlUdUxhQ/f
+agBRz8XtYpchYdl1RXNlcInjFaqaFPhkAXh5EGIFJBwNGt/UIR7S4R7ixRDJUJ5dwO/RMB60TvS
LKa16w4xxlhoEKqHoEbR7LolE4zgvc73lj3D7Bu3O1IwfWLX7EKzb3Y6/pjj22t3hZQrdRo9Ub5g
42PVTIX30qG30YLN7b/1kXJGRt3VYwRqioAuH6exl6a46LsDYXA/HM3zRDvplz5ssC3EArDZuRTm
NHEgcQfLrqvWJCHOUNhewt7fan2J77m2rUgF6l/n0yAMioWoaLBUEITnpgzT5bMwXQewSgy/sQdB
ttPLLx/cikepWXPXJmWGdzmU8qOGnx/x62hQgNHrnKnbSh9U1VS5GxafQM0WYpI1IA7x8v+P0aHn
GZ6uMFijrt93QjnfOsH8c5tSaJLDjmVbmzK5aWWKgFdfRDI3SvLCLCQ/iHm/zklxjk0FyXlBU7Ep
Ja9/yyrM3mtRHblVwE/dPOTNyocJyFMPPOaetE2nwGFKkA7jRb889cQHygEfK6H5Xu7lBLo17wbi
dvVTXt6DN8mi8h7IB6JjNoQJqf5qBD8Zr8kClRo9BdpaoWgVKewrk6JrBGC9ECGUKSgee0cY2jT/
9Y3+QdaGYNIzO92n+eTW8tHmSN0nqC5pnREh4q48HYZKXsrr56K5hQk6pgt6aIfKD2ZrrIlUEqkz
7a/W0dhAaPyZbQXum0/YYxYkecLa1GXx5gX4pukBeaoSGHxYh9FiMRFSyh0XStaRMC689AOKWehr
xeXhlZbq91LDQNyj8BanriWgICGfIH/VxyKAAYvfGAMA0IrtcB14/bEUOq6kX+lBlsZHDmKpSVi9
Ec+S5azuJ/YmsGdN1Stv60A/3vkjDFUFf7fR5wAGaAGVDIO9SpbbOqWvOFaznD45qu64RqcOruVj
zBvrMSSQkS6Z+gGCE6PW48oc9SDpj7GUWbKM3GdkQkYUtm3a5fUEm07uD409Ljj8Y5ZQs+9agvR8
v6OqOryQZUFdyd5HWWCu22xJzDn+N2TvR7GiEK+/UvmNHo0soM9WrT1TYVQ04rEumvWmsQaJrhea
yzJPU3LOONz40XaLCrs9A3kB3iMg9sYEj63BpQlFnfqNfqhqRBXxLZHxRk2QmMslCiyOcx5WEgGb
zRE5m6sXA1HCqo3sVNKO/62w+0h3/Wov6tamhu9uYv8Y3Du/a4UmdtUavItJ596dJOzxTdxG1kHE
HBQ48QIN/IM1FcyZmvEGDsEXlLgXeb2XAR4kkzRXwwBucUfwX5uYfsvlCuLgzmsYqVTBSgtqPrhr
/I8jUYIKsetLoAEN3w4bcygZlncU7MPeApWWGxt/iDxkI90a1E6fhw4DE4+dYzqZpK3spqK+qIYe
SmJtWR9PO7CNPLA8qSjDl/GvdOtNZ3QNJJds1kcrEaeCpiolaB0XVzKwVcwgn6flXB0ca6sjZB1N
xhJdN7lZsO5JUQzVmsTyHkJGEYna+ib0BSiLIQ0k0CiCowDulX7EVMiANNIXCgQ96lgAoTHT8p1t
SdhANK4ptNhaN6mpfUtZXrUlFkOcetazzja6PrHrX9boKBtvvYUL40LzZIeg0LqpFlvQdsy4FBHb
9mBPOCnEumleh28m9llifoHkBSkX7j76xMzr5ZZb3LvdXEV4VhJlbc1/EdniLJ9Lr9oa5X2FTSc8
HfOnDOrMMJelcgRGTKbVHkflTzJLO3SOxv+/8sFfX2LJx6Lp5IohsNycb7tiKAORfn3Xw9t1cm+Y
6ILIRGckvfjD5S1ihWfbz7INAe+8i4yJPTXf8g0yqWnVxOgHZSYPsUwBWgY6WCjlz+Q3dnPaIs2z
J/Vn4SIIJEXPsCIj5axc/aGs6kyIo+7ueyJ6KLtAVFslLf1V1xHIlLNy33/fNMwpM6ZNxZFELrpk
Ep0ewpKfUZEjokZXRLCwSwzbeaJecv9ALh1HHHsa688/RUde8C1eYzx05rwS1q35l/H1EwFRgwrX
Fxqxqf+MhdJHel1glTfZ2MvirJ4X3aI3erxWapsMV3SHu7MkAHMFNe6XpAWU3I/9P9mHbO/B3iq0
/jzA05jO3n3wHyv+inEEurZX/JIRaJUjFEB5IX6a4IVosaDqgvzaNxNVYpCYQwS5ZwFgcqf3/uoC
JHR0HRwd7Uo1xMrca6hgrEWHKx94+9HXAzJG76CUqeklfoRg39KOlfQrqDL077HWjDPhQzGwJLk/
fYhxpAqTvqBY8MYDPwMlaXLDK2eyI0tbPY5naG2QOR5cvCiIboDhXSgSUc5nSzuH3QxpwKmoD5aj
nltOuOb+Y1To0N8aPtjFW0eyicmF6V6E4r9YAQ5qeSSDdD9g0EdmO+Xx+AynTlhjhwzSTsptrAtr
D0NFlvuKjN59knIZWOmQuscHEyEI01loEg/pXrkDXPrWjtihjhgHOczpfMIlnNDAhd07406d/Gge
YQuB6beXYfN7JAl8BtVlxNVg6Nv48rWVuNFK0JuVcUOxwsC0k2iiUzf7usBfR+cBiis+GNLIJUTE
WFl3X6ml5Xk9Wh9n0W2Ecw73YuOQ8no5s7N8Rq0vuSRRa4vOyIjHtPTKNZ3NCS4tNXpfJSavIPxu
j5tJMVizMbr3Ds62yIwIIzh1QlOfmmP2+XlhZvQaH0nnIitBsNAvXD6qNasbsWZyWQ1ZN2niw/JB
m/pyguGEBFJEJHnmPWm1N/J5MLwRxpcZO7KYMz20Pm7qukdfKvmAZiCvp+8atd6LWeHf/ghUN/ty
n5mEaPKAz8afkCA3TXPEqGA3YsnFXPha5v6uBj/JdZ6wteheFXmFBWpheqFqwjs/1O6cQV7VbQk7
s8LiJ5CIe269hPrHfqDpG1Re0CZHxECyshHAFnTmMMl73bFQFtBS/w1Hkjxj1LgSVvRu8XtX3dHF
t5h+CIR5b0Y++Ebd/r7XhzfIWrbd38i1g52ZWs8Q/87GELNedc81G9N7Yh8T73CFnppci+ixr9hW
NRpTBhK98tzKMpHwlSMTmizvELpppRUVrqGNBgsv00NYvNVg/pnuNoUQYNwc4ZH0gMsui6i5vIa6
MWq1Sw+qaXWwvFC3MNANLzieUrvblMEOvWFaQD3neKtIsC4QOzbv7+7IcNXnCAKzKbmcNb2krEe7
RtlIJpYIfjjh2TKfmpHTs+SvxGhE/7yHU1+V+aL3yN2/WoUF+ZhA4qUqprzJcXijWkzDWtknIABc
YwB+L6JXYbFHQe7a/U2Gk5Xc01vcuj51Pc2pflKIXwSFtdH+k9fZG0GPLZZknpIkfo31xHIigsE3
MtdkPm1I1TyiEZvjej2EAOKSDjljKHSB8L8frU/QmmRbh38NrvnX9/wHls9iHpfmx9kqnBs8j0Ah
cQXJueYwq0AKE81oWrETgk4ZOK+1iFJTqDW4RibpwptAQoa6RZVHHA64sVG53eC+YDX0CyFU3L6i
b/qDnybfui8XL1DwzoI38aqChgtJRLJxH8vymMOrLlCOwq3nx2cOSWzrwwP7CxEQi8YLqel7cgP9
8esZgEcizCfQlYH8wk3Kg7KNzpdRKX5qaMwYaJe/6g94mhrTAEC6ljaRfA+6InCWBxmTM/8wFAJk
vuxKr9sPD+mEDJ84xsdh3AoOfHwEpNSMjI7gpqtoFGRTR3nRYRk7H3gCmMCGItNNzjo31/y6ilV6
cNhdKQ87TXw/qF7RHRTrtLmIcCFZqAdlU1fpc4WIWClkgO716G8v9GLRC+kko76WgeaUrZ9w4czb
gjItICV/UmITvgAI9wVgOtb6AY8EtlrddnpuVe6G/ncv3kjt9Xf5CvnkGD1/zIhsxlqw/dolblHy
KgSWvhVKxu2hYI4EArmEApsnTSTrPpy+/1la7H2Ca5KRjIIZ3X9rScT7XYZkDSktW6qq+J6navcH
jMupoE8Cl/GKY+bDGF7IknC9EXJJtWhd0AF8ALGqUjXkzet3sXpW8PM2Zsv6zsxFG6cTRkiK60e3
qYqB50iiHhzG33lMIUdruJlY1N7rn8L1q7sX6wnInb3x34YqIf2h2RB/sPo58D0bwg4goD0Fi15x
1g8QOjvhW70vn4YJj1EfMPWonW9lFhjMvGPZhJ14J2Kv20FOcbRlATUxKhiTU7X9wq2nRYjmpWvu
VETPo48zintknFN43RnEjE4lGFabI7MG5nNm5DaZTHC7DPRAJ7ctrzHOZp/mKke+pAKJZXp/W5Pb
lHJAcOmLX+j2gwFEVAYfrtJvPKz41C2CNoezaJ1DFyHBlkEDn/F/T4GF2N6I9sDwJ9FUlj/MNUQ4
b1gFRFiwtKHC51+7fXU992wSTnNmkdroIUk1jYR+fM62OcpdMHt4mGhY8AtRSKT8Ez1FP7nOxYO5
ZKD+jgiqMVlTlVfX9CobS7CJbiF+qN17oN54fTQttDkV4uF/BZ+2wbGuMl5cRB2DRF2wLXfDbIBQ
z/GwxYAZPYXr5vvYr9MkcJi6jQakPQdRGG4bXSUObbuFfOAdLQrlFwNnLOdkZntV4bsl9eKhoIc/
vbEbW62Vf1wVZ5jggxdeQBY8/0kOI0i3t9n6npLZcWTrv/QvKCtp0zvYKCcpTRSdQP+aPBfkS+05
KmsrDJaK+hLnoLMTPDmhGIt5RF0zxVTxIPDJkl1oO/BdhaW66EFUXTdyEK8NEGBlFJh2NbJ1gDbW
VAeb72M7ce79SMNYtGKpmBqiDl2lGyEpcvCnAKu0yZreeV2gqXo94l7nNMklpjh7Qr+FG8jeHyd6
6TMoGzKW5//HdsbZ0pM7ayTFl69NehyNEB4HM4P+/5H9AMWKhaSrHfcevSTINP+AfzYvnRFwzm8N
sEgB+mHxDOLwAlECWnUga/JGFbCOnuyWrai152ZC4vpY4TQKRuSTEBbIyznKFwty72Q3rORnV2p4
0oOcc6AU/FCqkgVKRAGroyW/Dw1m4DIXIIGk23iS4LW4B/6u8Eya67Twayp/8U149LczR+iVI4dc
0P37mRekMXJZ5+DjxlJk/66FLITaAihNI2KHwYSTPeKGQCykSWzEPNyaNQMEtby8+hAMD+RrmCbD
woUEmUkhgjTAz8wMkpIIAsDD/dfQJpPRujZxbglIN7mt60ivYfmsFSRSkd+Q5UVpLPbTn+jJJYIK
edoD7kUpRckPdeHUqs5Pz+fK5yD7BC0WbmHMbpfu90Bpad042HCAyudh9Vf8eQU9yA/SjFcqWleF
gBddKEcSOW/XzmBprB82Ay1yvm5IMDxVCMfgPDAtTBMpMLFxRtkL6sQ6St0ESDCblTxnMklfQp6T
z51mcJouGyk/FOpK7tEXDJxMNM7yJw7dzhUmO6Dqno2GZccNaKQy9iFJG0k7c1SGc79Y4bgdOl2P
B09sxWKgJx0u/eDFjGU69+e8hmZFsY7XG9wUZ/S1CZ0XGt/deu9a6IZzhDDapXHO0PRmR70YPj+a
Kft6XZ4/l/Q3i6lWr4BYgW6M/MtGuR7FRTRpCuBqIh/wMMnaec3vbn4hKyi+8RyykErZCBI8SlDq
RiCcy2D5dVuWh3rnBoW7IQqbDBWjmL/TNVD5t2G+TMs69TIglTZ0h0P1hfKOYrXhoEibaBjw6zf/
uEYWbVkT/zaqbCtHFH67Dfu9rkBs7Tw2LNsV3Yc90ddP0mbXdJXm0+HWxxoTF9SLeSMH6xwpy1rV
y68TCTP42/uApYtGPET+F/RBBQacyRJEqeRK6r0w/+Mt5nN91+N1bgbY644626zS+Eo79P9UK/ZP
Gv/YY+3dyb8p1zwC8q+ru36vG5iafyWgGEr3kvJRt8j8VEJXXI46ZOKsQciW+leEzqkgXEP2Aj+z
O2wjUcBowXjPWUSrLKsmgKSe7j1nd91Eh5iwnXizekShohCsHIqsktxRDLhAqjB4hoLP0oeMgreK
4cypHZMq/FibvjF2OZr4FZRmtOuTJm967+dZTkfzs8aS9dmBm3APXXsFjSsjfDUY/NpRbHxsG4cQ
ber6wuw4ziU9APhT34OvHiUQxuDNmdV32iIO05OM22zSO9Av0FwW3yCRhDvLxxGZeDJIZdldFHt6
PqL0Vnso2jv5dlO1U3GkV7CWMnOV7dRbp16FCAOQVkcE7Px4jP1nYu6VOTuaLXHtc5JCzViJDETF
dq8O8oPXDtkYSl1AHEOa1/+k3fNvSWGzd9uNZA+Bm7PixGmw2ALBaqY/0Iu3JdJnPXQnYWK9NJif
7XuTHhqxY/ml/zeFr4o4PxL95f/PDvH+emFYc5gx/hMj1YbPWrKUjzMiD8pgOGdQIA46RFndKs5E
m6ovBc01H0pf5LxnDiHfk3AaFCJufb5Bz/QX5jyXiUm+Tk5ob9OW8l6WL7kOFMyeCFWY04wJZ7/S
GdvVOg2BnsBCBZyGocFEA6ZrDT7Jy7AuUriIaNKaOR3bWAITSHuC6wRGoiQjULWAYIDBm3sWaxee
LaijbD+aDstKZA2vrzRdz9FMHXITtWq15YDZv1spjf24F6G+zVJzpa6XioR6rxPmnvEPc2QTCqtT
DJzCcsBWSJyjs2TpYxCjLKh0PlycjwTLhVDes2avNp6Y1Z6SR6BAkauraN52gLAuCbI9R0vgeDKq
ftND0h85dTcqL9/diP3zjAN4sAdKHc+BMlo+KAwRuxsJQauldhvqQZj1XJ66GnrXV4a+0EB+ouXA
vVOm40zr4gL09S6IkGIEpWKdmSkQGKS2PPkhAm6QHAG2Vl0bpGCZ5S14MAZRe6p5UdDuXgUpECm+
Sk9v+jZErNLkj1ChxVK2gVY4pNnh7NlsSblTzj5dlaefjonWIR8MIEHneGJoD2kAjfKCYV3GV50x
+Yx+XuSvGyrzOTw+MjWh6USw8o995PjUQHDhCKXX34MVHk8VypaEdZ/l1h6DXCB40ryfwAV/vFA+
k8G5WGUqBzTadU9E62BALw1VtL85Iv2wCbIKgGsbf+nw/CB6cRQ/rUzI7UtPyW0oJMNmeN3LAjYo
RWd4B3RWuz2Wr8kMcP+mNYp/o6s2gdmLIsbS3ihDbJpi0bL4E+o5+XDjeqM3+ZAzazq+6qpOtIQn
DcESWYXEBZnSdgaqmgOBCFR/k3p4UpiQqlMUur5tGf6nkfkdioZN5xaa2dR2WHapRmhlOVfOnfCm
5lq/bmng7BYxDOvxRiNUQmG2Q2iRqpiq+X/PqMGS7OVQ72DEgHhu5k6RfP0rHBitTtVr7g8lRE6o
LjDjnqbkpteGVHYN3kmlLdkz/oKVobzefQlFs1JJrOpBlwH1d2nXktdv5SUCziPabPOlm9nJvWea
Bi+NBX/Q6UvuGmmsyMfHPAJniTkcDmqlg4U3pL1UVbakJ/18Exmn3gKoa4RnMBLoG6WlpwiBr1jW
V7zQ/0bpm4zhvDWnSl9iB3l8w7/sh1wwW2l9Bs8PzVXvkK+MMfleeC0DPVIuzgyOJAWmOzdWCOw6
vXa8A4ruzEddhsr2GZrwEAqUSNCcp7awc7gaFOcx6sxhgK/AhL6mnerFL8ScEhCuBNmeWddDFAC3
IB1zd8utWIb3p78fxsoEKqQaH7DxMtMhVd0e/DCtrbHCC5lAaxE6MiyY7hPApdRGZERZx4FJu3iC
HKso/maX6Hj9rsZArbBZMmbfu6DHgkd4FSqiXypuZL+NvlhxyBUx6CFxOG0kmkhpbOEzHyxbTKjn
0rMpRsVf7ftINIdIc5fnapaDtp+OGjt5bMztXX5XbVt8Z5aa4USsgEJhB+7cWMCACt7RuJR8CYs2
7B0m79FhuJ6+vJVs+d/jyWVirQBvpmeO/vSuwKuNRUOvD1YcVMDtgZOW0LN9JKYBoNyXQ6zzlUoD
9OQClXZV7D1dE14Hg9HtJa+/Z1A2PzhB48g8sGupvSKfz9XRANJjRn74bJuC8ELcQEUd18Dog252
zIE9+LORtE5wt3E7saiXM+GYE7AXhWQD83L/eDjUujR6jFVt4KDP76lB0wsJ6mCVV+hMW9T2hPnJ
sdnNJfTL1iyGq4Y8DrujGtYLtIeZ8eKv+xqkPpAWXEdRJFAENt8g+Eo5TZYUNS3tUtYbrUqiuyqj
SQlr0Vd9Vtqub2hTQGswc7SUwI+avU45rJeTzaBxDhp0jnpW8gH2nvuxw2oqvbGpqqtCSSrjqNx4
qHLTWfaRJKNVPtEGAu8JJ0/GJu8wn/vTKTZQMzzsf5BZouBv/ooT3TrTJclv0QTGbD/uZd6BELiK
AvLWyVD0O+lQ4quhC5FyDP7t0joap+tfotzi/ncxADZvT2cHz5v9PJYLK8zakMQemCDgg5jIevoz
apbr7GoFjAz0SyJly7ZWKaWz1SHwmYQxSJ0iuTG5PTpTiUnQ17QMbvz061C2UA45GaYQHXQrkyKD
mK+FUDwHononlSwitviQ/TJ7ySEQZ9Dh7FsOU//eoSeBt+8VbM+tP2GtsUXKf6YQm+FNxbqbh3KB
CMGkek2cXn1FLaPA69ViTE2TsQ7rLJ3D9w7x4We/++gV0MoZ4Loi55IfP6XEzw2qjB+ea+c25A0m
FtP8Q546TaazI3jRQatuo7aesFPMvMWcbY9QqQyVwD3ud1yh82gbLcxipiw37LK7jjJQbGNhSrnf
NMzW7k8DQT6lp6q0ZxU/XUMTbM+wWezkZJCKpEtwRFJSs0NjwYDfkVtnQojvRqNDye4BQGYwt736
2qqvaUE03GSkksxMDIjDky8YxDuzLZcgEDI2AW5hVWh+JH4/rPODFXqoKU0/8UQXbF2aeJTbVL1j
EWJabDaeUReKlhfd3KGMuQxyQdqNmBW2MrMGLqIPN5IyyS4MRyfDRjxTjhS+OkvcpM1IZGLGxIv5
pNHjmt/lf0jdMYayKdVaxctG4Hp1hQAGLWZ0SJW7liC++19oD07t+tpLujSLbFGnLtDXCgf2SuSX
KV2l3sS+jqDsySjNbhArds0ItaHOusehlcQtHLNdX8VPG06rTxOXF2ylr8acvKh71PvNpON35XFy
c1RZHhJnd7UqJAw3qkni1dX0v+91S8sbyGae7vWUTuvjxATUPS9NS0dEiRr78VX5iBt/lZnv0+SO
86Qydd0ysDsqNURUpTnjmqkzM6ipLNDp0rG6rYVic9/0CsKJtilSeAk5pGDmtGpRlP0PMSgMuacq
905XvwjvqAKI6oDjUDVhYLfGSdadrnrhWQv0IsCxjsTU6QKMPAJKSJ3FoUqLR6ggpDVj6X+NmFHm
FOhAISvb6XDJY/RAfSuzMYWDMjZlBkHhI80/7TJCEh2Wqo6HTaVSVvbrcO/fQqCwKl49zIP/lZK2
wYVHvjbyv6rgrVqtdh1SseDWgSJfsS044NILfiKrFTD7SuWdLMGbdCT82L7vqXo9/IapbWvTFlOh
ExNHZYRuv4dEgvG5Z3VdcuzS4Lv0A+4xYDmT9zSGEoaa6GPuIzMg7WAY7wst33U7mHHN7/hSKilH
cNWvXAp5l+oq/PBcapFl7PNhIUhTsnwrMtTBPB/XrxVjIbSoUYKJ4V9NVqvhT8id5iUCbRPNZECX
Ectd44KPGgsz8lWqEJFeGCAufx3xB0pKsSR26FEnv2FTnZ3Vbe6ypk59/1i/XB+iQ5dMD+ZAb1vO
UJc61Mmw1uRTm8b5aNoVhDxcYl0RyHcFRKGFiaTYV3w22H6lrio1xy+FyKn30dl4CVrc+JNuLcpc
LoxFFncRaBwIpyxGYHkB1stahaAuM1YEUL0146z83n+Mr/lH9PMcqQTGRIzpvAFnt00kyrUZmG+D
sOJvKMFWt9uR/Y7qgwqByN5dUXTfs3JRywjTWeNDcjBFNI+BydFMGMp3no3OS5nQbuRWYIXL4UHl
3eaQ16N6f9Anl+YqFV5FLpida9rg9wc+f28xj295pwksgPt1c5RNCn9BUyqViVKwSwplJok70j6G
SHar8T3ZXZWwxImumGVlQeHdk+o3KKVQIajwilPZ0kdGzr8X3YD77FM8AeEAbi2qL+X4oVHesCmF
2kciP+WbEe4JGRIFhrXZAkiuXKGYo3iAzdlYAT4ZI7k5dzf3lczJZnQzVQLMuIiAzBx57X76M0Va
QB0uFof7ev3iP5QPeI+NFCkOX5iSJ2JpHjTtMT2ollCu2GW0Hm7CYH4yBaXYd4w7CCmii2CH+2X2
UWR7aInwRIYuPTFn355pzNd44JO2qIh1eaAFaN6PmERhEF+yVLTfgZKxAAOC7GQ3/MNwWEwMenx3
aKlwGmG8g/Z8QW35vmdU8aaf/5Wc4BkThFCwv0s+eFZ35zwWN2Ujy+W1+xgG1NZLq1Ezog5OEaWX
f7HQe61uB/XIKgx3nlhesGH+L3cdwfydp1LT9qMimkkdare8+z/EJ3BJ9Pzb01f/1iqKkE1y3thd
Fi8Rk/uFwo2xbQDbRIvS9Kc6v2TyrvZ2Y4oTOEo009n3vOWcfpbJk6rag2DOEf8gox/MAjcL4v+S
byvKKCiFqHV1Ec/z7+/u0BBnXW5iAdhnYp6yAR2zn0DGijqy+3Ob4UIxDMsx8EswnT+cxBPVd9zr
uZQLB2I2tx4rjvBi3/Qt8JudyYO4F9/xlkR78xxgleBUYEGzYPPG1cxKXyMROFxw/z04LzgDigYt
Z1RNQRbSwrY9xxLXdUiBNdc7EDgPZbQiqwVHH87/dh7Hj3+dqRrMtFe2hfdYWFZHRcNgTwx5umh5
ADFpwd4oUnpFTmDXrkzuAzdTOiw9tTZROJH+Jy2cUx0gRP9065Efc3OmYRtaEPWcHXh/+5S17jFv
pQmnLFVJ8xhelEoZ89uG91+VCLmA569CViDhrkvH7SgRtjs0hcRv4aXUokRL8JaDD/9xLaYcvhUH
MnNpwPyQ0P4pmKKan0MHwW3poaTwCYI6wUU/VfZxP6abrfZyGABTXuLXVyxuTTgrACC0sdVSpKFL
HzYo3cpNA8LiceLIZZYDYn6OHHvi9otcafb15eTbAr+1srZZ+p66rdPiONSar3w3uG1C/dF94LUx
+m2TPB6vfvpWwJluQpdvEbUfCUjdNrfMI4YYQKb3yIj/L959vaNua2Ebv0xoDs3YKIjTpSoPyu76
pvFx++pugNitrdUyOxkSyl5sYfiOKy+d+3/+Pmmb+9snCXNk3+5FnNsC9ic2Y4UlSWXuCQE/hEO0
/IAChGtWYElc3gyVMGy+O2oPNXfOLo5Z0m0T8jk67epY0+8JuIzD/F801pbu3lQbOvW6P79kmEeL
5Idgb79LuZWPncpoUk3pdIuWpOIlK7q+gmEizsDlfDOaMGxfwBdh+ZtkX0/LYIYOAMBvl0LgsED9
luiTU7e1RDkI79u0846QF6I+YJcvtCsLUUsZOzDrA9olHUsdSh4K1I00on6LG/LdESdGQtZiBy7x
O05cuqSIkVAB6xd7vmqpxlOoJWxJ9XQxQSvweQhO9c3hCVoj+y8AICy6/hoyjzlrIAcJaTMDxzDP
6kIdaUZs6kLzNftepRRvqDziu73eyQLnvhN0fYFWEroCKmMTRekGZZxJpDYVjmimG5JeJQ6lahtD
1Ba8M+AmuDaxseVCj4W/tC6FZ/YJKAawjGmOeEB6Hud20K6eFnhrKLiqUHWp4/kQA0hTkGqX65Ih
QqsjLBY8BsXow1T+d1ZuGIjk/QV751yb01cs5yo+Qc4qVqGylQVJpWgXbVa+2vYUD+UHjrKIT5z6
a6XYkL2D8sq5hYL1ZVIU9nkf9kedgbYryhJTYtNiYDiu8Hg17pKYKPSb3/pjDN4+sNADWssTfHpl
E2fn+d6YoShttJW6rboIpBZ6M8CF/lkr4sS3ENF2SSi/LMCYiT8Uq1S9kryu6AMMFCKST+Fz+dEd
7QlCXmrX6HGUSLYYYP4nG/tGZuKLwF2draJ5l6QxAOjkWn4jGaTtY5E/57L08DCuSosFnHCpcJr1
HNT0HeSJkcgQIvhmA78ksvJLIIKN+vXya2jxPOe21q8MW2BcbWmzPUwHBdb6xPGPX0q1hVPQFazI
3MiIu5K0pYJ7MvRf2BpmbZXzQwa9rMfeF2/EYPRiTmD2aXTyH66fLwrP0LuLGgQhmEprpMO+fvSz
XTQv5TdBjacq+zp6Df7qJvwNsQsKxfZ2Gz79YeCPat1sH32tpN3FidyXTp+fxcF+8fFxthSfRwY0
STJgJrYj0oI8ZBZUOet6bnAdB46v9TCltV7ikdFHEkDOTWXDCxm0Fg1qoS3wg6hFfzuEEWzCtkWY
YCPBOO1UMW1ZZwYNsriX6X+LW++Sx+YeFNERtQ5FBtnbnvIhQc7YAoLuOSeG23Y9VMiTSzERG5Ey
n7pmGcrru641q2RkeXRQgqD1SiJEiKR5HjwWvKxlqtekGa609EgPg8rko4EJ1RUdx7w2cjOqpG31
8a95ZItRMQTinmc+bn+ovQ2SKZf6PhF6mLxLQHqFaZy1YAqJXm8aEvfYbRYcX7/8osKFxYawsVZq
gJESM1DBetVULjNvKr17Hl5nt2KQNCcZkzKypjUaFYxBrnzUB8bMDX2Kx9BqOYLxrGJA55iaa1gh
kXOPrKcMTZTffZi+QPWNqhpetWCa96gV1Uutp08PoOeO/nGHT98fHETcCNd3oLO0dYC3z0PXDwum
kTyPaLpeZ/nU5X1vdGCrT5Zim2bT2IkoEW0QKiYN9EZ41nwCP7P4bwF3KULc7DkQu9fryvW0u3gc
w5bWR3pxyD/cQxOf9KXrkVBUbx7+4ZNfBLSPJEEC2u/sy/X4YVrgrBfIOlY=
`protect end_protected
