-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Uo95fralpLjXfuG0CZkao/ST71oC5/dWksho32QuF7dzRHQCCGMWRtFdIgU/lGm0jSKY9Ul1yIx2
PzfGun9M3XNFvlbNDngSAHwRYQq2WRg6/YrAXkvVnvShtM4u3w7hw4kTcF/oYmZGsFM2LzN8CV+P
lpowK29ZILPL6EM7HKPKMoUwVR55VE98UwQBxff8li/RNoluw9TnOWEXy52bD0sA6HJ1Gt+PL6GM
CH++MH+yTuElXyb9qsG1S3zPCY5hv3NsvnvTdZPirL4t3nh+unYaMfdEYx+Yk5OCAFa8GlzOHUf9
MUusul7rP59ZeCBfQ5q8R97A5jtDUP2oXPbxEQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 25264)
`protect data_block
EIylKBx/HwhSlSq/Z1gXiZjXJD+iWQZRvUCZ3vSCJo2/mNKZnyKrLbppzZP8Y1KZAkPnhxmPuLe+
k6Z7icd7Jf3lFGHFAa/fqcLpFpyYWOKujqxrCeXDmXEZmZTLRyD6IEMyFH68TqKyY7w6tskgjRDy
0Cl6tVLPSpe+eNWTcTT+39EoOZOQV0BL0F2IEYC0PnEZ6mQE70bXPQhys4dUwjDcDMkHBICYvnpT
x+gkkRPechHIEz5jSEph5HihpHGdxetBsYEKn+8Ti9oX5GhDOQfcOYUtBz9QtWqUKVxlIUI4IUjh
AD6NvLM7m+Rkb+ku3HkNS+whEmsIYRkfQMKNwftXwkzNzlBHOXTYt7kNU29viHM5TansIevHbbTI
S4CMwEiu6CIF0B2tTwWOHw83mMgNNLdnT6TcLp8WH+f4O6ISWcAl14fOzc9ZNbOdH1Va8xi+YlJh
uG2zgt70BVOuBKVB8dyLhLui8Z+/GzWruMVUdKF9qHyTxoePJYaCFN8kO0++jAelOjXcOVgd3y6X
BZ9BL5E65LB4YFLSLuo5bRCY/ZiiYXnnTQWwwmJpYv9hSrTbYTpkZx8DB0Nc290DeMMEGEOWBie+
ZNQBDq/pxRsv6mHE/12lDzeRSGyy4SK4eWiMykjvchHEzInBZ8NnHHngfJypr6HsUuQlRzcJ0yLA
l3ADvoIOqGCvY28Vudb6TBK90uRYD6qYp9ZuPM3+5RS9v2GVMQv6HCPPyHjanHXO5ZKg9demckNB
qfO6BXUy1Via6CaGJne82Q6NE0900OtuodE0DLOIoIbG5RoXzsxTkXvA7C0LQeqTvkozvYtwxXy1
6Jgr92i4UHk585xvHqL59VvwafwygEaQsbUYf/ivhilAnyqgM9Fe6vLecF1FedK6s3UyIPi7cN+W
WGpNYLiIRkYs5APb2hcf79w/i4EqV1etFE2RYkTMlm38E81oRrkWCHhxKePi/wCwY4uIU3KoErbb
gXE+g+Y/Is7YxC5Dh2RRbtdSA9oV8Xjhn5wlSrlkQbu68Ifb+bPA1RVKCihjRDWft2fd3prADte/
mhbWDnynJ0cZcD6yLOATWhiEG2+vrZgSqkT54lnoKINcv9/pX4sUnSKDy/TUbdtyICL8oPhLFCuK
xX0fnTTXgsdIj2K4AzzhmCWikH68MEnmkqp1BiPZvDNdaQfViUCNZkw9E+D5TTqdPQWY7WjAfVQP
ZaLW1DK+5aHCijl3GW6ShEL/EYFszzB8Lf3pyqE14FxkwfEP+2KmChmEEMaPFAb+w1m0dcFjtpg1
1H/Dh2qDs8oFPsZV3EVHqWVpxgKx5gdVHB8RDYCI2n4zgIDnYjxxP97Fu/1Y2wKvSLBEZ+Q03cI7
97QATUchzPHkG8/rukhQT9+3PbAh46VgpOglSGiX8DA4g5Ex7JAlznFd+JfcvpNh8MUb5Hrv4R5r
bcWeiuFzqLaWXoHSBGO73bbmmqMWMm57/cFuTo5iC0phKgfw7pD+wMZZoU9IxR9gS0lTY516EErm
HQ/WQSX8nDD8WpU85DZQqocFNsxbtlEUnSUUpbw2oBm9mcB4NXz05/VrAhttsIccwN8vP3x9F0n7
akL6g1TBwV64niqVfJuCNQEL7XKZeLYi5KvTDy/1ftQDmwBDjTrOTOoOdovh0nwHG4ZDDRLYBEM3
8HmnX0jJUz2cORmnJ4A7n/vCf+0MS8Dt8K5CGV2f50B06RG5+AYnxvTeNSqInUY0QkjWuD5bNWnu
slwt65mlXoHdtknp67rz+WdliZVppa5Yo0LBwD/nTGqggChZDEqh5zlU22rY8NwYd3kSYqNE/eq2
aW75rePZ5QQGe0Jaf5Mc3XpYMz+dLtNkUhXbAIXZFhChHb5k74It3H3WJhaVkYIYQI/+u9zWAbA+
qOVsC3xxn51arlu4rB5yUNebTvf4Hvy92CgjVpyOZAEqr8u9JnRURYo1nnXEm9ADnos4mYYc4c+g
XbYYudAAa6b+WWwe75f7NX6A8oz0MH1dO7TVYV2yFN6gjKZWCpGcp/rhH87/VxMXp/i89PV4hMNf
zARwlcYlAusAH+UMRaM4LbBnhcFLW6Vm31g+SWzNn9PM7bSw5sPsEyf3dHw8Pcq6ySgL84bb+wqT
xERO6zZyYG/rBQeF1z94I1FGjHL8zkbSDJJjQCMEab5iSXuVFH47hJ6VKDiDGwxE86a9eaoJZObF
HXK6W85xUOEdUhW8QP9gVnlyR0rIhLJ34Kb6LHDDA/DRSFI6isxeEyf7irRBPCou4UEFPCYdVGP+
zEdydgQGH0F8P6ADSPRUezvRPJbWjFEjnFo8Ko4S5YEBvrCXakbopC/V1un63O85DVfGvZJBF43K
0V3lLcw360XAW7RwB8cISvaLUyxLxoLdlc24UjWI66uMULTl7OAGmwRm8TyHO91S38cdM3gjjRR0
l9g3ehZvCclgpXEsFirM3RMOW5KKy1y4cRdfhaW8OkibrCu5HJFNHK40Aa54zpsDhB3ZEeP1q8tb
2xnyDR63QFV6GccgHZ0vm/t2LPDKZ4lDSGzsAsxR5Cyuo1t5h8fH8m7XpwSz6XNx0G0ZPYcA4pCV
U81u2Lo7WO4Rrtu/pl6hDOyov8qhRCh+KnosocnbYDxhohAOx7DB8jQh+zAv1cinklCSDwJRbnxh
igGOMO2hjNhHOyR4vl064CCpdxx2UALXA+sXN+2t7hMbaKP0YUzHsfwS0UPSDWVbG9V23TtlqN2g
HzuYj4vCuXzkszqHEQwjdinLWZhkWpIQQAG9ydkHNvyKjiTkr0W4ahQTLCZqXneE537M2pLUXyLE
+9CDVbc68FDp2Yzsc/p31NW0k5UI+lit31GrB0dunvC16Hl1p75miFmndXV1gEy7qzx2Me9eQaGB
R0lfRJwZxyRwG5PweZZogq/1uoAE6BODcN8DTAWRc06kZteGEAGyO6X6Hm2hp2UF8BX2S3kp8c5A
tZo3vqs5PyoNFSwGb+q3RRDPHJVoa3cS1QDQzYy7Vba5BH9fubDKtslkRRAzZc/lVfWxykMqR9mx
eb29Y9ddgqBKhwKPf56XO1rMf5JFx6YggJxKaTBxlAVWq3auqse+zFm84XW/jGls70Gy/nMRq9RA
+tC0hScVm0tkk1FWPnKSI74nPgZbxZqugMuPKkjmaB6xwqFilVh9cEXYjQTB+1XBIwdqDp4fFHFU
H9ROltgTUz/sbxCseflqnrx5jvwN+DZxthy8sO+qjq8BdlwrEoimD9tCjteSdewIluXxEdJA4LAo
GqY7Szq/NPgrdOVVwq3swFEz4pUY+24b7kyzKnLAbibB8GtfWBS7T/QW58uODKY9gB1WOVKaapls
rYeTYVMlJv8n3Si9LPIuz35yjcyYsy487E58chuWBXa1SProl8xLh/QWB1pZLW1CJFKn3J6oV23k
bU8GWSSwqQSa531U+CF++tIDhctw5L4Xt2uBBUo9ppm2qSfgJq/h/NscM8mxInSmzvaH9Ohn2lvI
KPFHdSipzyYH8jrgl+XFUS1fC5ulVh6liFaz39IDd/eHpts2uQhuwZSYNU3xZdTQA2VeNsw+amol
lmI/dwVtBqL4hHw9YYWqfDlP14PyZxBE+QRdoT6PNZveSleu2OUMlEUFDT9d6YnDu1dmpMP56BAX
OYyLNzwUtidB2duluEyLi4VVpyk+bi5+A3sT5tV+L+noZ+l7/jC64CyyF8JYuZknCuGnDofJ+BIn
GVJFSGfU94ovbabRrRi0MiYTvw5hBuikTuF1Iql4Zqv5aafSYK6MhM/UGPW2S191ohBX/8GGFC97
bdH5yazk0EOTrBwLMPANlCfcBDLlsrPKYyY5QwbKuaDQAqdObV5PxXCMykGlxsF8Ypu9AxYDSnRF
KOjEPk2cmZpHhByYYwTJnbX2oNgaw/HHv0ZnUFNGBwGL9HBUQp1Xrh2K6AmzBDufC6At5d8TKPdo
vXLqBOddQNa/s+qYfVgRdn7BCuEu8fnRZypHOnOW/S9tyzI4MFvHMZHTUT4mzUBEm0RNwbPVePG3
7AoPbaVJfo8OOvFX/ZFiVZcNDyZxOqLMvl/fqYMFxh46/02H2WBtPZXTbV/q8ZjgYCOpyu560Nn+
Utkwgr8buaVSO5Usr+ngTqNegY73OMvD5tOtC/BA8mRdOE/olRHD4bo6NpLhysiWGK73smOLeSUz
+KBSv+zsr5qIQiFVZLoWr1u7Pz+sxmBvWEZl53BEN7oa7T6prTthpHoKmZmlRhAdWrCqv8+anHA+
xSnEFwbjvCoBXJ4qhkKszBufVhGrY7/zTVnEJ664sLETvGtzev7YJaQbzC3b5eQPzQbgQxckZbk/
0BgyeDIjUPAchV+FZ5dppn+oeiGmmwB2MmL6Avu9OUEtVd3+51UduCYJbSZuTgcMOrYX+nmLQLkJ
SBPmVpiI3oFoyfijybP8sYkOHi9jGqyjTcCC/FU3p/S56io8Q3fD55sFPD41zjRgkcE6Gt1l+Zfp
ouCONZ1kWnxF8UWSUXvrXf4Lk1+TUH5JN58a197DKiCrMifOK0breqPVGWKih7c5W8j67DvZr1Qx
ZGxe6T5Nh6xgdPUjf7tnbpyiFU5K43T1tUR9bqbvg8EgX0AiqWyKqbouPLg+1VNzdBa1lYDFLQI/
iYQdJjQ9DmXxPu+Rdq58YYUTrJPglyV2c4AuEqQUH0Ze7wvgFz1p7DtbLifvu0LD75RhKtaEZKjz
HmYKBNVQfT5rkNG9Fso3IlfRgN+GphmKhFdyTJDt2ie2i9XmM8bXMWAne7/KeCZk2Cq2Mxn69nAP
mDr+GxNkFbAyTMGEg4+w0uTUXZ6rx2cdaWeGk1+5V/6rySA1AmOVI8Y6UfvMqJFHiYyjbAuU/iv+
UmEgnmYvwECDRBSTEMnZVghFOZ+yqiH1wC0SFDYT9OVhjCwxmrOVBJK9uRFrTH6lNQLgC6dUmnO5
6Ef2rbEGMhYz9vSEyzlfgdXPGaXJzaz6fKlsMAoz85j+99MI6d+xcRfGa3rg2yG8YqXX/WU+q19I
FUtn3ol6rcZQXrmv/lCAjPBbCsE43yXrA7Girm3mvNRyy/g/kHx9PsX8GrdUud2pgLXukLvnGDK6
VPU/qnoVmghq44RqORND4WtfskwCsNnxd0TdthXKIIWBhXllV8WdVpTacwDC+BlHM0oUoO2lyv+n
3KaDCXv/COGW4RF38eZQug7fXaUBymjOVy9UDxqbXTCpHx6nM2w4fcw6ENcVb/lN/QDb6RhAb/ot
ACI6DSt+bv8vmKMY+vrlYa2hGMrzZ9NPZnRB8Sf0uW1uvmWbrR4jyaOCTpWh8ZYQU36ZG9l98zyy
j6eECZa9D44xDbst7qc9xSXdGmkde/oRlQb80qge546LBGLRcHefhfIP+zr68HJ7/ZY/58yTiY/7
Ejr0hH4AQ42N3jaZXOIluyvsvq0X0Hm9Rz0/inkpKtjD//aJ2oLbHmfwWKTFBFyYYivlNQlEPQLr
EiGB2XIm12uEFej2WcdWRlme9fyMxHh2b9rVwxK2lglDXBvKw02BuYc4/MATgmp69QAa3r2HGHZ2
R2WEX1uhZfF2yoc6gMA395XBJgjy6AN3uD5hmnS6NqDfyRkAXMk77jxltj9QSFJa0Vlkck3GDxV8
KjedofRwRXhpUsYlb/dYlo5wXvkdvt3w+o0L42rt0HFp3etjd4QLDnKTTmgUZemBdCqH1ab4ngiZ
MSReuQpdx9i0fq8ZSxMIPYS1VGRDRKbtcww6iytvdbOI2hM1WgsolumbsLExA7NQcslW4zsb/Jin
3RMy5UXIZv1tcq6IG/Rmmd9wS9HrSMFAf38sliY4TmK0zTGHGEw5RihGDj59xuNlhWfQXXyTBtKo
P/mt+y5toLGHAlyuVKdJP9Cjw7DkyP3/vJJ9CL8imOuMPFZo2Xo0oA9LxWGPJC50vfNi4LllvfP0
YsrcsWsjlVAC5XlW+CapJDLiAeGK03C89yZg0PxYCGHEe0LSy/+O3S0p6PUW7lsZsmHLhi9xWDEc
Gpjw03v4qlt7urIsJ9uMgtwiC0uFQpYvP5nBeebdHUmt433kpOcpFoIBXCQjsjariRkWP5sYUb9G
pSPWLqMsYQCbmecheBqwtMfGgg8g26fnHPzNpn11ymelwPgfeVxHJnJ4EzjtkMkMCFKIoGdTpj4d
sQKys1mrxWBEULmcjGkqPy9hM5SElN/O0eid9db0MWam1afHh5DZDiULFKp1+ziU+1TT8hKNcXoW
QhkFe2kL5iYhM+ZGbZs7xfYL9aNyVOheUKV9dgMmugybr4XzBrOyXJquPzSPtQ10462fc9SdP6yb
bdGB50m5vHDSDnwwpI9kn5AbXAG1GIPg2EjmjU6p5LNMChQkxtQ7RrfeBEiok1yypC29TtM6u1sO
b9JCkIb4EpLH5JSkOPklLEoIDE/98cKtfwNCGb7dk60pW5eQ5tcxkDMWmyBdrrCXGEZIS9jitDRs
6OxzhqdkK2EqSSySBx52bB3FRFJIM0y557yYtHIxw77dz97YPpL6Yhq1P8MrPo4wwxE9y0isKgO4
XTQqQgetvmSqG1Ze/38wzIb7Mvk1Kfan79GBy76LpHA/3cRtnGl5qbwTkfQM4kQ5CffXlP5TvV3R
+soZk+N0+uIAwqKV+23/mIl3v58yxI7M0o47dAsL6dL1yv1E5Irn5n/c65ArhsHf98Vdme7jv+2n
zCp/Te0xLp77woy+KybMeRLmjxD10yAHospWGTkCWB9F04SV4d3luRYHQM70sOLMlGcMwavC1Vmw
8RT7t+t4kSrv15MinnN/3yJwakClymO+TP0EAnu8TFyGcLAkWGcuaUDl9EjWgJWl5B9K1/rVZHZN
lTK2O7PgJUCp0L7fWE1JJI0U6pEYgAhR/ueJjcmgvTwwyiL3M5HL9V9ENf8/Jxc/LdqoxjLdxO6U
m2Wto8OrABzCJQ/IuaMKldVeQopMIv1D4DA9w5UJrw5Sil+VeaR1n6//sir3aMSMHt+OUT1Lu+qQ
e9BEt0NvZAZxUDBDH1TCoqXzafrXDMSxZSprAHo2XmV9xv8RG92us9VAZALiOIwa7cWbGvg4v2sL
Hsqdq6lTrW6VhzF8GN9bcvjtAtq3U2+hGBG+lLAmTxC1o6Qw7QZZeYSIv+zWayQEl0sgchVjS+rP
dYokSyLido6fpzcOIqrQtLVGMzZLps61Hew90S3r+EfVPY5+ARVUEypicTjr1DEzdK+Iwlu4xEj8
vtKLTZfb6dHPYjn7Zql0kCWZtCYGeL4q2JSeaE+NvLFkRVfoxAayNFVLCRBCh44jtcBLJU5MV7/r
aO83E9VR3gqMih0Nt+9RNw2aZmbHvYwmGQWiz0/Plb1+vjg8SaNrgW2vRhBZTFhvhwnwXy56zHJG
I7d4uHJwnfVfW/ycVkNkJ+/yF8xwtD+HxxC8jVCl6ZNHrLXy146igCmOElmLIp15sxztTl43Fwos
4TOUKUT/jGMWJCj7q4e+UB2YqZIa5Ao8Sfs9s4Wm3EFFRbr6isCKC+bMeoCMqA7U3qPl2gv0uLjV
GiF6ateFjJ7nLwefgpD9km1u9GOX/opvmDF2o0IJBMh+U78BHUblNxd+Tfr/ktKqUw3EKfi+geH4
a2gof8AWox3VpYtfceW6Uoihp0h//NxeBbXv3nlSYbFMk0X9XyCo8O7LOrz3UlZWydYs4BTerhxl
Yvggxt2qOrFjLF5dW1Sf5PKrXA07m1nnIP7WiXssb6ftwHjsaj2yEn9yJX5NuyQKoYEed9xiESaZ
5hgdWet1eB0f97jufUqwM/eBHaTKnZR8DxHJvb2uHN/XfBkmjFiE9lTL8ynAKPq5L/2heSc2MBZF
RbnTdOzeV1hhxzqYrxo+vVe6e2u6oavu/3lMr+IXPMi2fmTMUx4XnxNac5qGbD0E6SKLmoxbOpjd
W8IExJordJ2uqGJKCbW/O0EF96TXHgFXYZMImc6o6X7E/rpgsNKtdN/q18GoMoyhpvz00QRVTUz/
K5WDo7amJaPv2xLBqACgmBbqndylFoCD8JQ4XUQ4j1j0aecsOgPkpjp7d2gkEMrUime8pu6WTDcJ
4TLoeFRf6gZI3bjROAjFwEnDLRFIS/rlgkyW06SIV394/kUARAdEi8W/ps+Dji7Uo1Qika8CbeWk
/3EJnqS33v5AiKuFUdGSXfcpUaUyez87kfhos+hmDsxQDpqCdMhoNYaUPS86HuazzSur2I9FWMfl
4IYwRE1C+jyLujI5mP6ZvMwLF7E7bftIZ+zoMSNQXh0QjjjN+MbXdxx/y65FjdjpyMeLKU1M9cYg
rkNtG8E3Oj16rjGyqmJnF8oCtyiXB19b105ZwaE6UcEryCCA4hi3zlBm77x7X7wxlC8rpA4fJ8Qs
J0U4OROl+pU+YSpyFEwDfaP8Tgb86PKb4WrhI6dCvWGG5TU9xOdsNkMjBPtrQu+BmsY42vaNrusn
T6Dt569WvEJuHzfOcfQosMcVMAbwgVWnEGi560bC2lTAirMsQ6o2LQZW/Jeun0wMeNk6hhkx/8kF
HuihOcFYr2RBC8ok3iXdhnu8TYLrsL0QPFo8ID/LZIDd5UwQ4w4w9Dk3UGJi61RBwxIAoRpnufrr
YYpleaRi+IUgVL8n/IgjuFnba4Cz9eNVY1OI0Uhu2Qb+aeHKQxupykwjHPxh8ML9kdXDhR+YI5nO
9sq5RF19xfVGwtReYoL2vd83lNJuwb8xBEqW2W6rCBpnUBQki0m9GamjuVSOBKbtiUs/c6SxkXvT
l9KXd6k+lscDanjtvLKa007Zu5g/2if1U1ukH1e4F5t6wGZrqtR0sCh3pT7VLmUuyBJwpLSTBISD
tvFeo9Adfvr78sVoZ+wQBxvz4Xea/EMaIvuGBM17oNn999uOiHbHjIOCVJinEL4MQrqKRcM3YB9I
FI5DAjFoO1L+ByRPQcYOBhwU1L+WMXFn25C1Z4ocVusesH4IoJFPT76zUK7Wv69wlNeRgCgUWCPF
pvU0HI7tVox1NBQaatBDVwUn+lxSU5hjaTG5c8FgfrmF/TjUWy1lsuM8UMk5HCZgGTtDbSo4wTF8
kjgPbjIeahbNWNFZLt06TO2kFUJQHbX4SEHQb6q2I5kzUMKJByU70ZdOeFwxVz8ObhxmSoG6t34r
3r5dR+SMGJasbtAGJv2s8frxCltRnULFGKbOgKsCiBXoYz3ge+7K94LjnMf7ueARIJexscZvguUi
4EeC+79JwsqzPkawPYilAT9eZFQCARRfJTVYHolkw+XkQLe7KXuVTEu3mLQUYbWhdRAuLB0UrvO+
OHI6WCSFaH/14fPuun4OMMKQdnFq/rnSA9qztwSbFZdqXGBBMbk6bt8w1ISgMyJh7PNqyJYgl6Z9
jWhsn7YFg/Ddr9rSzHWs0XNgd2doZu9zm0um1AEdQwVczkMg8BdBR5ZrRV4aw039ImmvK1WJ7+Li
xNLhGpmnBIQfz68/5kPH/0GeElnbRgXbsEKrpoCI0OGU+L387tTQEKOJuVEiTrldnF3is7Nfe8Cp
AntopubyIKaRTxrcQEPECMKdytmk1MK5eXzA5Mb6bMUhrADdNyF7do8VE05hnlWMYpYNP/38APeq
UQng3vX6v9i6G3Ii2bLsBIHfbEHYhwuYxOfKiCjxduB2pTjcYBkVf6hCdg4M/zEpkSXWlgGrt2AH
3NiXAs+5GGQlnl4/mMIPd9yKM0PWRulamfObbtXhvY+2+JBkhbVi/yVNpctzgs2e9jZQZeuFKmJZ
VnOmAZqe+ufdBxnf93BZCC5FFMTvE6hkviw1lm29T2H9ofCgLqlCi0VocTmXkgY09l8WR+wxri/x
mSSp2daHkDxomw6LUJyJJA4vEIIIttYvdJ1G3L7jGyOlIZlq1G5qfJvBf0BiJ0AsWqWnOhRvVfhh
wzoNVq8cx1+JAVDtF6/BgMeuDecJswwNTQJ6EK61SF5DWizLJP0bYkhYHvQ1GG3S/vD7/8k3U8Tn
S58yUkD4kDZZiNomDe1OW57a3Tr+IQY4pfT+Apn46AJwZYLbZhIhf3RUu+CWmzMtAcexGo3FmfcY
kVw/ucI+Vv66tiAWcE1JbrR3Dkz1cZEjuv1Sct9oML4rOEA8WygalBq1USzxdtJHkx6A0rpXzTBP
ccTRgGVz7TCQEt9flkdJhyZiUo8eK2+dPMLXfA1xnNEL/ZmD5htonGuhY5OicU5CkQehdOOdbFVu
MGw2iUrvtCFCSp1eTUmDDpjjTBazTqyZldeGl35mtkv0BNtQ7MYxBBoZ4u+eJoN3BlrlZWxiYnLL
JWZkg4ivoWzRAkjENTimnqqDAXvyQdCHCfNcGRW/3sL8Rnrpixug8ZHpwLEOslog0CGWcNtTFWWA
bXYhIpsca99+v7JeywvwkUO+Ukcy0vI89oU0HztNU6ZiDcbq5iNxaqoNyod0KoPks0z1cmSg1SFf
FCrLuUEtffO2ANff1zdM4QcIAtrogNXOjwDvqcgPTaCEaAuNlDYm49/y9KRZr46tvlgMxkPFmo5J
Us5NAvRlemFMCb2LX1Db6rRo1mewN9KlJBLLfoBG/id0eung3+2v47sjHP5dpUMaWG8Po/Bitqim
cPtf7xOc7maqKDjdsSB3cZpNnQoF9cmsFrJdB9zJ5d/V/3Dotvb59nlNAloLSaZbuSrcvGTan2yP
MnUbvfdokWIs01V4vNHcdcavMMUdE0Jda0tCqcH42J/3tuh7A61p2sRrofv6dHx5N5ic7iCZD9MC
Zwh1UjJ/d+Iettdf40c8G4Gx0idp1HxGh3Hcw4PFpyyrFpbVM24UXUQgyN/8eC5yYYq/xKi0GLas
lG62SXojcTu+p4OSpfYAHgE1ucqQrQOMJZf1PqOCUHm85VUC86IeUlpU2LbjaYH2i3xr3AMnC8/o
UpqFa35sjA1e8lEGrI7+1joIlGn4ta/aKhh0uoB8r1ghYTpqT+gghkFACjIH2nA0vk4ZUgSIALl4
BZg1TYJvtW+G4YmA34wKAjqBYTWurqfJPQYHiEC45sA/Nsk3FjsqjvYRBHw2ZI1FSCClJN5CgRZV
nHRAcejPCPMQ/OeCjoLlvxZEAijzktGMJv+iKz1jUpaKtf+7OaX1+nnxAGFYHKavszuHpgITpKmI
1NXv+PknJ0ewpfghxUidBRmIE4zqiA48rwikw8NQP+NEMPtSOk6+q3QKyiUYbC/ViJQbWPc22Ie0
Ri2RHy3GtKELAIYzSgRC3K7j2C0GS6dWU/IZRmHiOEnGA9ZvX/fTq96Ffe8cK7O6h+DNcsLYZvdL
vL8O6PhrIorlMX28CevkX8X9LrID2tiqNMraUMHf/EhkhLglCl1mJdgzvb+08k9XxWoYECd2YOEa
dCCLfjol6E+r6aG1BfYWgL8DtqMJa1PWJZHhNslyZI/My6g4/tWLaRfbpCVZmOenRWHvWAjGss9M
OzVsmGTWHund/vRaM6X2I5ftW2+JtAdE5MGEMqOeGxw0DJ5iazBtNxgU1EQkCxhytpIrUidCo+ED
AJ1YcyFG2T/6Q9AsdZ2uQ9wf/NNapNC366fBzem2WAZQS/AgqcQ/6YOn0XWtyRH27+BUnooQ8ygC
xzzbBge6Lso1Y8GmD4tUmGl7NhlWNADxV623gmOi4QmKUPn4otuVNDqyY45sbUGqeG9EnR4d431Q
o8cdniDQ71m5Qg7imjUyURqBPy1cr9z4a8dSB6BCMFPJbNr93OVUb0SUK8h1yaPSEOWIcyy1xqRY
C3yhYGIzh4ggvBvGcrjArejxt4jQZKrJdwYlRSiju4FMPnBF2TcLV+7U1eVVUWrJ4pTyLM4R9tYF
MFOol35k/bI5+RI3VSMrcEqMRzrEFB4G0Gi2KXFeXjzZgHVdhvYl2c3O7vilsdepuqc3WA5jvAn3
vW5mPkHLEkBQ7Br+Ay1kLOCX9BpkfzoPeSW3idAO7fUVLZbMsyr4Qntvk/QB34Sx/Aq5sgV80ww9
qbAcMzMqvJ8wWqJhuTrdK9ACtSeyRkv/GslKcqph0XX3A+WTa4AeP1eyTQ/qmb8o+jtUNjiYEbfh
AK4QcumJ1nyXsyFETPVi4CMjPkx7hLbkHTwtXgnJ/3OghJs728MEaKOpiBUtrdE/rk52CEFSRyW5
YDnzcfTn1vNL4eoiy+hbOWNH+qFxk7RY0G9KsxNROvg1W1UB7FgpF0vcOwzh5tDjZ7gOhAeHF1xx
nqiT9GnDBWXa0m5ZH5b2s4q54OG0HVx1AnJ5EdsperslHbGMPvN6gdWRXuyi+l/8Dz43qKKQYUBV
VGmhAw1Nbbnr2twW87Ofr989Fn+gfte46SsNlg8sW+6dpQb/VSsxVvLcHnMbPeQ+cxDPFGvnXYQr
xitwaa3Jq27wsbhQo5jaufCbHZu5UxOtK8STetCDRAADdNVgTkynLAYTJlT+UmUCehUfYIDradhB
YGUpvjUNetgv6xhsPcW6uL5yA4T7R+Y5L+B/XoOz+rp73gfGwLrNzsSsfSsftylsuuGWhFdi9KuP
/NmD373LAaX0cgWUe3l+xkUWnBgM/rsqkumcX79NXSGqW+g5W7TIGyrm0+KAZxSnN2Ts06x2hYHc
Kt4CG0qV6qv/yyXraRmI6eE9ff85cg1b52qXkHf/xcK/b56HSzeObqRpIeqkkjkPbntn9nFZPlVm
MNghXYcR8EkqCJno0BlfkAzjD4hTp6Domd+eea/NgkZ12i+KSPRYUTfRAQbEVEJFwCY5Qx4iOOm1
WeGMkCGVdwJ7w1ZyTkTe2HlkjCK829RYIkODzpxLaSe8gqXX5ockVYp54h2YOMQ4tDuCd5h7GY8i
3c5hpt0N2k3eItOvCSFGEbU+InHpK2kAvYaJnXSLYzD1BKUqrBtyBKnaAFjzzCD0g/wPnam99Ym1
vO9MSMr/fQkB7+G3wInmErjU1y9DJyNyrEMya1riZ8hs7SlIXauWY0PjjClSe5CVcYkrPQyT+1cX
vHbTj6YjPFqcHa5It5sgsYEYEIGENHXmoIJueLxjyYqtI9W7Kb5MjVW2jMCRZKKCDkTEiQfJH5GN
aPS4PAZZxTnCwq4vJEInuKZtaSwRH9DXMvN48WDAyWGoh52aYpe65Ku+z49qR+z/eeUVdo9r7GvF
kFdqVI99x3F+qfMJwQyn3ogtXkekD1C9qr24igs1nHJXpyBqZBkbHaJWRWOvcpOkcE67TLAamqSl
yjHTl6ih85aa7vstEmA20gKR5jpCOVY6JEFQEXvHSvYvA2N4qNJ7DRIcsS0AeB1oygSdtLb5xAMq
WGX3RMP0yCw6DoS9dPwLOx9DH+CK0ht0422Eews2B01uB/qjhfQE+hOWHKYje6geEHKSsiqjx4sq
P7G0urpR2sHvcRIV31cqBykf/HyEtn2FTDdtSWsCp0NZyTUDhuqj+bU+oSxgKwAdV+5HzT9Rpb8v
iFc7r2KgaRiPJPMcv3qiiIh8s3ZSHRO2/mk42yQeGZsObPX+VAdM8TgAXmKbuya75kTlYJzcwB0f
QBVUtRKXH5T2iJnP3JZemEFenH1FKloZXmtkl8s8faAC8DwYmeQS/uBgoJVaMqBALKSeo3ZVEYTo
sJc573dmwXVzFT2BBAD5Md8eO3bdzrVHqHe7xdXzY8wdNhUyIexpmGnVVuJH1RfK8DxCR0CJJCc/
6wn0U4kSnGb8nLuPOADvN05JbXAa77FTxn7wO2ImNQKHHFDKjuhPOhfoEqr/YTxhYYy4CNOZF5pL
9N+shtpIJW2EYxp3k7Ub7jqeqpxED7TFd7lRkzi6v5heIvgMfdttJiVZ2Db893kIGdRD4MYQva/V
oiJNNbDST5ReF7fsPTTY+/V5iVOa01JMrV7eBy451OVBWRAOwoqKl1O0DgpqtZ067eO5mdRk1khJ
23NSbn8NwahtVb05l7E4Pu4/q4avUnrPTIeE2qaX/KoFpnoWsd7RV7HRBzAkkSlFzgJTMA6f362P
MJ1qm8dyHsPV2s3VK+EwFANuIEnprE5QBsI5906QnXN9TsF2L7AEVqEyJu1ryv31bOS0lC2n47u2
bmkYRY0iGbHfQ5EAWDQc/aMVfnSZnEizR5llzw7i/QlEBtb3nHyZ3DWnYU81/UTFtVWuoII9OiVj
/D3sW+9NLBhiUReWDjNpVKIF4aelr/0WnFuZmrBuy3QsB5reWsqTlcnQJGaaA+LKcblBwWp1ByY0
OmVc/zj30JCfsWBhQAE6AvfMFvglTwCXisFz1VvM/ToSzQqvvkhWB34igPJ4n0KlrUaCjmA1N6i1
YOIUc2VbHg/4620hpQsCRxrCTqiNdMxDByIDVShel/trCgKh8A2N01deUZnZihrRe3fSDXrB/ZBs
lwffQaVHVsOhRHJurdw0dAvjTsyc+Y7WNaBRtQhymg4RG2niyVHUxU4iXX43eLQwwF7SiCAAh/px
I6wK5m53PjF8DejctAGVDnjUhjGQsT6WtxyZNagCp0jW1SHiNNnDErFT/ucV5A4GR9V1ejW0x8qN
ZbNf0Mz/zDht5dhxgdKgjAic5995LDT1KSXnTyD+mL+yJzVYc3bcqwq6hKZq3ETOi+9YA4U/q7Rn
SymJakMJPHteJGzYi+JgN1SZs2+LVY5WqMUDX5qYBuOip1BclWe4iPmJmrG4GN6HlAuHKwRoIijZ
D8g92BTu4h8b0eHBF9ZIUc2KjtdKx3OfnVwkHoWmSmpZDmA+dngPcBzykjMg1SD6IkBzrw3gW0A/
v0oFFANTMfZpMwncapW+IDFmrh9r26yKVZ64AWvf4lGkoEmq696sCgJbXZW24ATteq2nI4L+x9pt
yCjzgYmZhi2kMqztqID3S70iOOFgYga+GJGIGv+CSQq7LWahlFRJkbQFuKKCOpoeqgvy1kI0L+EW
4BMHaOCX+1PjLDGJ/SA5wB9SGoMacM6/n1pwDgpXpmXCjO6S5IHn+/WH31nlaA2iFnLcF5MXzKKj
pa2qst68svUq62cd1oY2KWNUBckLq9YtPU4BF2ucpdBIOAPswHCSc+1clIRyKx4ycTqP7f6LO10P
fhlGTRS6dz12nczX7Qd2lo182gMolAmB6xK3mzmn8uKUZyFV0mdNAQIIqR1QDr0ci8/eDA772H4T
Nel4s+RfprhvoWXivLDv4KsVnAo80uGpX3yyEKd55MEWZNH0uGAJh9GB1J+UuJl5QoXO5/m6niwe
mMClRc6JHXsabjzpJhIc6ETJCp+mnQZCaTlqjHNJnLkExXJBsIJOXBuY8J0Qym5CNOkF/W27oqyR
JZKkIvQzKntWVtOdiHCuVTRbcpcfQY2yKqMszIJ4knSZL4pZfaqhe76DKWSbyR9M82MVpUjNEjQc
2vUOjxJVwlm3Sfu6aguy8MowU7o2c0rB+S2xUdFHi0BreDKQn99sa0ZIPFlVh7bUxvJWFyjKCAE2
wF4H2ZiHI0sM0Z5FtkeyhN9h8KQQyUzbx2LGcbtX3ExAsi8RUnkLkRL1jma0EZgmWgwzvcVcGCI3
3o6bfEmFXWcQj2pxlCEJSgB/gmxdIWwrIbT2yUFRgRDayTPxbXyd9ARlpvHKpJL/yC25f0ERmdTu
O6iFL0BcUhw7GIxsU/hWqE1yAyu7kwaasg9vh+WyZclfRN5g2/Ssd4XKrjSUioL6V32n5WIzyuv4
rq1+cmZRe7uuWCOd8ZljUu7edEm5pUSThuXzD/NvoA7PowvrS4Cb6aVDNJYtFvlL1hTAYMQWOvuh
qHzQjDHXW9ApfnViKGP26erUp3dZgrjJpx+fOlreh5umjbS1JPDmatJj0vIEkNkUpM5YEsqbb+7H
W9taxB5prl3XRb7kZBg3uaKr0ELYSTqurGfj8FyjnZKan65Ett2AgMFt6+Y5Leaf1DJ1/KydZijs
bnnWZMg0gVm7wIPZY9t8maar4rffmm0i4O+epzb82eOpx74Bq8BwNZfSNnP4C0x5u3cosrfKp8g3
TlAHio+zxiF3GgvVWiPK88LpM9ffuH7Jl0vPbV9k7GGOrPu2LhvdJesoVeMD95A030FA4c5lS7gu
rga0QvMM0cob/3tyLxXobvqoCVrmEw+eli9Rl9Wa3VBwOVa2xGGBTD1MlTzzyBktnBwFHNTqJiiU
T+0XvEywbyh8+kEleoJpZMfu7MgfANjZuxRoL9hjB4bBRgaIz9j6pYTtSIVDSm1WgiVnW7zT9jD9
q+KVvH1TIaehGr97CRBZlqNJsm/yirVHiMrhcagfgXn56cFidsQ5hRVEn08nSl9Vmvh4oDlYv2B5
DArwnBskprhZl9c45RTmfqDXE38Ck/oq3ggE/8ZB7ZlpM2e8HpgedcPfNZeodbIlrlJ8gqEiRztM
TVbWcFcihN7ttMqPsyzbaLhl/KWYVQQp+xvsfkAxWvU4eLsvx4zxLWNtqlku4A0aS/PIsNjlLTqv
MYE344e4Q6nZ1CBMTGMGOuyCKkOOPmAR+dDkuf94TZqixyVFWsCHZeYxiLTrDY10ElrGuQ56ZTc6
H1zZASM1PEbcTKaf2zOP0N7IIjvFNbhNdicNVNgWL1nHtpveLgBv2X8Q2HvzRMziBJj78SmonJi7
wdAkjhPobTZ9OtWAWo4kXRcnJ+b3aqKO68WNlKTWdJXaMo4Ks2gu8CyOi0NNHbE51YzJb4ywuE2p
YSbNjaCRSNV+6lIowBw0Jn3mTDlpmg25MfTivuMrgaNuFGssYNkUj8UsBrWqyKSAwZPA7C4S94R2
MK8YqhWiOumaXOW6BZ4Bcu5nQaKdxJ0Q0b114xb04iO1/riguM+2Wz0szKTnxnOLgS8oZOi9CucS
+GbAo4g26ozF/9Z+dbiY1klL657rcROmxkY5QMcXRkVX0+AnsRUblzHDHsg3x40gFdYiHiXUnhjg
LvxjVu24imsnIP69pokBTISqBk7itDXKJCOSTaua9l3+j3wt5WArnifoaGnNSeHwOsEj6aArPvKZ
vJwyiOhFa7E4xnyMbDXZFK5a7aBKFx5Tw/fAMGUB2pNTTUix/eqPtPLBwcTxmwmpi5st1qES2qdh
Lj7VF/+LQRgDfw9CAqv/JV/nR3edpg7MCnAopOLjY4GNeTEOs01YxJdC1EiE1/cEL2zjPkHNYsew
h8kG0Smb4+8n9yll/cmT6GjHv/ItzcMTJVkaLmaFVEWhoXxzBCQD4VVurtKUewnRzLV3pfYTvsRE
6qsEMvQP7pGuNQqNBx2Kah+n7pFikFdu80jHM4iUyQ1XXkyhjaWJHcWoVshnYk5FBqErFqzCrWRd
zKb1Qaz+9+93oqUQ3XlqRrxiYq4txZ+IiXO/TJDc/5zwSpfMU0lz8+/jNke/s44K2Q1G0jEs1uh6
9aDGKW1ttMbC/+HHz05eGidPt5zSFhvVSIyjk6/QnMyUEAHc7vMPxEQjy7nLgkDztrUt+AK7d4t/
4I+AxXBLo/XOTG4R1hJl5/fWb0gAlCUC4kBsXpDSFmNGKePe6MbNsSmD5oGRNGn57qCj8dUkwi5y
hBf63CU4c0NyDGn3D6Xs1wxxuK3z7I+DWjsQy8isY+0FF90nwgT0xRwFXFuIOxf5PCQH7ixHtgRr
iUQQl26lRmuGLGYI9KGdRtZbg8b3b+Tg1WOkCrQm5c0cJDQ8cIbNmShydYjslQ9b/g5CUeQzNS04
vjw4M+OCHabts1nTit1rKRStbSEzfC3GyBYaaD3fNugjG9e+jeRHEih0nj/13Uk79SfR/sma537+
Jpuo5JASS+L6avZL69I8hpqwECUgeq3uuum8/bm2wQECddzsrs9rLl2tCZG+pFSt36Kad/hGVreQ
AZg9frEcXZUJzztKjZm/Ya7+SMN/oPmqwG18ftyic/WHl/I9GoWOSz5UKjeLbTXlqoJbir5Gkura
l4y7FhS8LnUbU/gSuAjn/Ke3rT8XjXXG6MSSp8JU7ZNBM0j/Vl0GIF08/55+HOBSR6W/nGPM4ORp
KRmEzSsOp9Zy2ElS9b1URlQDOPlnTq6mOib+BvAy1cWW9+hAkaJsoFSBI13WBsYHK8HxdNWeU9/X
ayZGGPKJsNEYHcry5EYkCh+c8r8soE724aiaHG80gVpQL/JXSA00CjlGXmWNuQD6Btjlsod74Iwj
tNBTA4RN8Lk3mkfLuSqNWPOQmy4BSY0R97Ag2/wrU4Xyk0iSJec6ZER+/C1xAMfY0zQruHCVMQvb
aLGCTHi8VtLBs9zEhZEoK4pFCNzU5lukhIpn3C7vdUBJ2Wp2rv/xuH/56MMzdQwecF7PNlD8ZNXV
QRyufo5KdcW6paajQ/c9Qd0gN58HLTK0zmFHOEUVvlBVx/MgL8NG8IjWwV+Rb0CbGs7/6j9V5uAq
7jYjEAmJM9CdbsCFfTv6IaatvB0AXAq91I0KdZN0vPR1pOAE1J0mx3dhlvzwr7d05cL41jYc6P5P
9MGUuffXS0yOuHAl/rPY55802zm/5n0xpzVXw7kAvx+pmb/reKL73NA/0KIh7qoI89Le4Bt9hTnz
BaSca5+ERsikaTPH23Ibg05L+xJWG7PdxSkEx793tuwFuXyo1eZrLzw20JWtQv7M6N9mvGCsHeGN
JOgykImfbU/HqMW3SZ3J8BzRkg6+8ZXToIF3DWXrzGLkE/cTeKtkaHgtua/W7NmCRV8s1BZ6Ojkl
7Fj1Lq2JO+1uBPxrsgDlOlfG3nWbtyYIfrNxpjpH9dZw5bjRhDfcB6ZE1jDRN/+J4emv7cgnHfz5
6bt9Kl0YkE8mEAa3yZ9l6Hh0KOqi5Nw3dgXMjmP93TftvhF9M2IZmZf/BTWZRRyLO25DgdGGmdx9
GSalIRniAUhnTeq3lJZ3ctiKMLsCtHLuN3p1DXfs4m0LQ7h+GNV3rABxKwY0OZoP+FnZ28FWJkFO
HK1veRE2DHV9fIBb8f/M8oEVdF69/uhFezISnYdknzZmBY/puOxLCQ7LMkYWiF7mMCHAAOrxERZ9
Q9wncsX4b3G5m8kerIgHGlWIXb9coIp33w9/HGtvA/IZp976fkaPmODeKSRN+Zom4LAt8DnFIhUg
2RnIIaJpsoUaqRTwWgIsVZE92s9clkmBz6gQWEUNk0fr7dlnFgKGYYTu9VBgJm7R9u59Sa439V34
M6W9P42vTXsq0VLvZFguncrK9mXfq2qW2q/adLMhYE+3dbHE1/JWPOeysgkzj4yLImb+svXzQLQj
tASXRXOg1Ek1Z8EXBf4YkHva5dQUPKfGfoJJY9Ql0BjaSNYlLkqcfUIoxi+8kEWk2u6+6he1FijR
J7fafwigm6y4xaZaR4pkMliVpo99zX/aPIHyj5VmzZe4JiXUqF4E2dyK6pgsJfOj+ZH9XoTJwgy6
r39Mo3mCAqsm3SiEuE8ZnztMJzZWf4zkwQweQLrWzNj+xoEiTKknbT4+2YJNAH6SLY3ZctvK1nlH
6RcGbGIi1ljYEKtvUypAIzOh1NpDGM8ILkrnsfygv1xrEAO5eK9Kx7NTLWFBdhuCIts52zFLIuVI
D3+I3H/JnK7XIz5Erc35VrRk2I+gvO0H6P+IvqMEGjhM42/kfQNhrKhXvSpqT9WoN+ePCz2I5Ncb
XKBlEqqHR/+tBUeWU1GfKQWSgH1ZsknMS6BXaRLz5WRkgKF4FwAa4y1dWNwa1YcWNNSlLUG7ObWG
n/bAgdtIKB5Daa+WjV7HsDillXvCs1FKphG2sNj/jO/aR4tSdmmRxPj66b8X+eZ5nrBnp7iK0TYK
lilUNilXuZUFwKyZLNqetNuGeGZ4RjHhb3hhBIZJrkpxj+pjnK/gfjChGl3dc/OkZEpGpHTbO78f
c4hgEJXJcWEQKP3GdM3pFLdx/nSEyGkvYtQa9nN6U6QjwldSrJHmVcG8gDdkvoe2qcicTpUAbC/2
v2ebDxs3+rQPXI8mLsRwfXfI3AIH1AZQJ1iQ89tDSlI+VPOD8dy/kpskmhLDLT3qn806EJ01+d3a
Psb2yyrD23yxEk3hkpQCxIj+Vm8zxT11tpTs6Xpl1iU7GESJdlpt1ULSFBw37efZC06cMIQ0nDUX
mB8tyN75oIhRLbtuv352vPhtbwsc93QeXs6QLBFnCpew7zsU9PjWaLuAh3/EAgwF/BJM61dwuSOF
K8DQbVl+yHGtM2I2eaZte2/ta6rl4UpBRTUAJwe5Yb28q3Tkti1Tv5CbSCbaf745eld1oIMc5Z8S
HY82s4NgQWJTAzuK937eBwZnHm8eqM3sf7rL+3K3ja9A6RNFvLpYhlF99tqxxnGQ5s/OEMs/Oo4T
v0YUDa8kwVsCJghWVXtBKZ1vmLg/x0stGKPeyqa+C0Dqj8b5NzRg6glBI3BtYJdpoe9MNAg6n7hk
6EDCsKojDEjtTl+T1BcFzaGvpfYpBSWbfxYOCyXWpsg/huDlL2xR4SJ9gHWG2KzXIh78fj4zxd9C
IvDOeQE8eDzIMOV96xN6rXGOVvgu2Vau+wSA7CS+6Vxrq5X4W7SfaxzuvV7Ts+JWCMidUVZhMvN8
DjFR+dsWv0stJfliafPp6HuYFCHqMNG6DqlM5DVPKmAmfs+q+OkeHRAbXtsMFDt2l0S3aZT2ifZe
CjSI0cdNo8RiZE036IGpfunw2EqERouYzS+kA63U2AdtHSKHkLR7ROgWg3xTlk45CBpNEHsZy2GH
gp957R53bX7dKKq/ceOpT59AsYBnTfvVpEhKoJWPMP/o2Of8zUJVY2krBhOQYFBerPLiyK1cNeVx
JdlleOHnmPe4xVTVSHLYXI7J1y5JMiiE+gVIfcjnUnvPAqT2si+f+HGV986jFvm8VlGliypsIjDk
ycv2jukk2v6vy5picPkE4MfU69KRfCz8fRpcRNHgYRlOACRZlvbGzXfnA2hgFRpDckB2gF4twOeh
umZa5oI5HMbEjPuRAe44h04WfwCgoTwjMdPzcUsKkg3v+01eJ397vs6ilZTesKy47LO5Y/rPOVCb
YKOzA6UhlZRed/+nHuP7ZEZQSLM1bkJf0S13lBBgDZJJDOuugOiecVGtq754D0CVJJDGaoKHMyMc
qaHn+dYPJj6AMH5iGr6cbDob7E2Uxkhqf5j2Eb1G1H0q0++x9S2kT1xq0LfRDQ/FmPES3M6ZZNcK
mgWzZxHOIistA4cUCxeZVmt2sbMOyiT7CwHto/Ok4G62b6Oit8np5X6/5/zKConRmX+g4FMIQ5Lx
fe5s1DfvuHiCRwmbNhUcPXKWYY0ORPHfDi52k1O0NcDWR+HgELfeHRYs2HiAfFREa3nBhPfMPRBn
LFgn+Tk726DIFQuKkyZFfbgae4iHC4krYWk7SM2SwFLrSLBLPyO7YODRaoP66X456+C0xA4zlMwb
BHQ9X5dbi1qO1JaO/j1e9F7ab4OQ83/j8tYmMNS8zQYGhd5l3uJaHhI9X3ITYnN50CBaZfO2m9wk
EHflWr690fnmZ503PV81LfBJehQMvRolcf0XUf3rKArvJwl00SPKXzdWuooPDPR3ZGrrZafEIBe0
QKS2vmt9mYJR77n7RuR7d6ZoOdd421h7kzENRiU9on6BVgXFG6uVm+GJVoIvD3zT6brX4isXWdBP
OdgnzJPOAoY9ux8R8d/x16CF4ZbL74Tx9qKhDzBpIscdGC5zaaUH8aGu3sOcqsDpxeo+L8ETeDIo
jILbRKoIroCkRcBH2oAe8P3WnfWjLfY99rnEx6QhNKgx3ph1KO5UB2igPfTyLTxNhnvYSSkiwEiZ
Aw/yUK1/sKTyQZiCVc3PJ475OPt+ssS9ulZkE92uaIvjeZhnUDR2mgB05lyfVwE2A8Vwtmll/8Wv
r6C+gPHUzoprjypzI6byhXs2fbR6Qh+CoAXK3iIz3Gq0HWhUNIj8Hn36fMdEB8Njmv0pJaVuJ3qR
VfgY7tttsPeVbw8GzBboU6mACWhbHtobAHEU2fjwVkhF/fBP/7YymUoef6UL1UFKqN/wZQ54wDN/
Kg1ZLrcd9+6LM94NBLz3YVMP90+nQjsHTijduRS8UU6snQhEwYRbcbeVFey3tvsRZk8tQR3ZHL+v
g9M9CGz6juioNIh+qAfe5bp/LI72HJJoxtPRfQz/BM1Nug/GLUAQx787xQD9D3qsvRmWaUbf1A+J
flKlfNMFGbIK3xBWWGjabYmAZyjH1P9GvOvBQgHYntwlfM1mlX3FlVAYLfA55bjDx8iYrILZZVMI
n4Ot3UhWtuO7sYclpacVvS9QLB8hswIQkiaAn3UWIYuiJvTF3qhQ8v4oGmARQSCOrIMELICglP2w
ukJ805GFmhwLYDMdCtk/XvCqxbF7krNq59xEd39sfs/jldanemtUHUfrQ8tRUmPfgnSZDNkpF6/d
tzLcPIdU76ryajc5DIsToIFSRcxWmNiWOIyRzEB5OJiQPf2thzi6IYmxAycQhecLgJSaVrSRA9B3
TyywI6XcrGCK//oocKeEIsA2ZVzFi/IQ0sIpbNul9xg4VptN4HM2HCmIHewBTPRdNZ5lvdNPDWAk
PFJQuAGsdJy0BipNcqh4goBooAPskkcMFitNexdlhIzs9D1fd+OThRk22Yf7SMsZf6YtufEnMHni
ynVxdzVxj9auv7+tc8ObUmFt95NNrHDBhz6ty+vzaMg+IzfwPgrGglwhuHpos+3znwzOkoBQZPzC
83rDrMHpHXYanBpdXkDLkullG3kLCxkygKS3LXdC+1IPt+5n/JH0kaNaCJNzxTT4EeDHjNr3yYEM
TSK6OWIFeQt2STV0Kw3q+4+/hsiJze3BJ7+CUgsgVAiaY804a4R25RxNe9yEGBBmpvRs9I92fvB/
8b5EtEmh0/XvEAxEtYJH5lHwLZi1tzjvC4W+xYsufyRrBVBdal47HE7qKg3+nn9bW+Fo4Gcy1P0J
WGfY+oXjdoyGFsDyb1HCELcoEjbWBu/zqioONcR6z9YGoiGxAaDYZIF3lghWOoA/l6+Y/cKfw9zo
0iGLsMmm+4LpxuzRhfMtwmEjBupjr747FZjT3lVySLA+/ZEKPUR5UCqlucUyOhglwQybpsLCDn+T
FJb72cyVS3KjgqpjvPK6IQCUsPvjWStSvreB373yJVTHZLQx7rwxkMu5I9EAuSeL/MPAM1yOKlCh
fMTw2pD21t2PiltKJFRD7F1PvdzbrTMk1K+PmdoIRWViLBk4Ntdnh3eJovbJnCen7PnxvFqCw40N
ySuhkveDC8rcXOLDZTh4NGLLtmPPNW08TO7HbTY7JM6QnqDOfBHbMv619a/AjfDwfi+AcGkBDzHj
VjFUagvz8jbWFr3Yqdn/xLbf5vFXn7GG1n3l1kJgTMpo/mlbUlfBx4Nx5pY/9yT5T+RaW0yJ/Oqp
dnfPrFXGLvRDIbR0WqavQ/OLyv4uNtxoX40nCEEJB4Ph0uSHiknFMw6S00iUQUmYjYVgsbo0UGs6
5Cu41cabezVYmSg5bq0zwzJokAu7jljQhf0s4ZitDap/qWogePnV9wl0lOVBpb+zDBpzM7gqxNBQ
R7PzF9WYsKLseRW8lkigLhHkohCEdJ5FFqr6VoZ4TEyQGG7GCpv809/13Fa/3sxWrU47+X3zgCzG
KSHJhiXa57g1u26266gYw4KF1CnQdvplO9xh+KKlMHPqHTxzsavZWYHeFTDffnEe4PPw43EMjhI1
LgDbj1JIIqHXcHh9XoBV2nFccqNjZa9D7MBuBPCfWYMbapZYL60h5PAuwrj2WP2CeODRPGA4+WY4
+xxHJ+phvBrH4LkqIDYcM1c62M+bqOfgWmjpdZcDXVZpJ0Ii5apMHzgOJVd/Iby8oY8LoJ/wnIsE
JYmtRkR9YqFMZigz7w7hmNXUfj2w64sPukMIaew3E55c2nbMz9ZSmeX8eYcvu1ozSAp29FMzvP/l
/CsQ7oUUZ+uHUAeZjlf/Y8Qc3ZaM1pxgc1aj09zajF42pY46bTA7VJF42UX6OG4qCjATKF/uH48H
J3qBPvSeR6pj0L9zcv5KpuX5g3Q35S7Discd8/TQf1GdzB7h8be77FX8chXKdVG1cczvLtEOZeoX
VqS/7w/dRV/SNGka6KoTfGHPxaiwB1Xig3BU0OFNPf9ukf2oKQQAx8t3DSlpWVyK7JCeXRpqGEOW
Pa0eF8NeP22QBh2iU2PMk6uLK5j0zbCU7gvY6uoTeyVc46qx7Tl4/LdMyhgonXcrZalcEo73WmoC
YAA0SmDOH47NdMjhgjq88AfZm9xsF2Lf0+GRVnldPsq3yOaROpmY4CPcXG5lBcenIISB9IAJQ/v7
2wS4oedaZ3StVAZ7fhSklMWlxuBzBPXs/3qSUpaAqh/VRLf7UuapCTxBLmrNqJzGWUmrxetTJuWK
fQpOfLDZCtOewfDkp4OjNThcSnPb4gPP6BtwgtvvtNcd5A/4WJgRja7w5sEf558njl91tNGN0nI0
bGL/v30WFnzRZMoNawfWqLRWjNlXnj/YwH8R9x9dVzUFklKBgo+UG7kGYwz9heERhvfLH5Rf0AmS
ZxgRFPxPBT8X9qhUgTtE4+MFgRgDqZ4mKLHxPGQGcY+lSDGoYaAHmlOBSoTD+dJi0iv6cm7xDxmN
mPyIw0PSKKsNPCvywsg2L9kr0WChlraCPhCeM5+4RDXAgjwDntLgXFAXwqmFSnWveWhMHrZaPKRp
Zu/SeUZkeNNqbaL1KN730uYBFgdrt2woBRfyK/b81UQhi+4jjyAN0/pnopJVZyBerTO6rA1sw6gZ
/6tasY1swff4ULk6d1i+yG3IOsc5ko4XwK5GLphmugisJXF9bwKyP9OsQH1IDCWH6JSkeTaxcfFt
iCE0bcnansy4XZmZgEIcnCmcUc0gRBX5ITU3Qq5wvky/DVRMGTrLXIQaX4qHU4C8noWXAegl/CC1
TcpndYu1DfvmdDCMlO/peytsIrNqEW6dU5gNivCH9HrJ27xi9/xXKaYzBBM1cfKul8s8+P0/eTHh
t5qEytqX55OpnOTEzGJqcItD2bYLt1d6KUYkehAhnOvjhu4sMx9TiCm79uILUvENHL7sSEW06IaA
2eGoqwcsuYLcPDW+ngS1QQGs6Ltw9Zr94MLlHNy10OdPMBneqIKyHokVDqnLYJIrdQ7LqGvXaH25
Z1p4riII71G5LW/uHJSDq+Lrd02OdSXFH4Ks9x7Cj8Z+p97iAQ4kvIhv+IKIq5hNckpZwIgctn96
lbrahjtLnkWLurJChKrVcjdoJ60VltTRo1VnmCqVnBDerZxXcNEhYLHOWiNUiN5QYfr/4jv3/nbG
MpxUHr/ZCY/mYY0sp2WaLXVr74BAD3XwU1s/mjvMXSoK7FY3+D7FY2N+zT/v8+nLtickDOg4rpcR
BE957wTHilJ9uyssw3oUiCaLydMFJVHYBvvMs8zYm+uodXt3Dd78h7g4P1A10r6c6uKimUuAkztZ
SuCOerNWGDvvTNbQ2HwPHx5quvRix8eyXEaAP7/XeG1z+ckK390AzlTXozuX8o2dRRWyoyBV5HQR
7ITwbNbBaJf5qjFZmepE/5tIQcSRPYOsKLL5Ba3mmTKANN9DEpok4/JUbopu83wWhUpe7pivzgpe
RPuQtk7BfjU3cEuxPv+2ZpRr5EfIdFXhoNYqVfppnf7M1bkKVe2SUCBE17efzlerVfVyK0T3gTlX
LQ/9BUOUmPupi1bC4pv8ju6bW1n25JIm4x3G1teRsTqQFPFB57cOcOgsj7g6G49jjVQxR80CpoDQ
iFtKwkZbWI2OEpvEtB6BUsNGqBo6+ISyzegYtjcoiN+yZMyt1ZdGE7uWCHjUx/qZ9KAX0/Dcmzh8
m3DAho5kt3YHnQIKEpyG4h5QcOVReBGKVkvWmq0H54r8Crd5RghyVeQO8YFbnNc/gV6yZp52yhiR
gyG4tfzI7Ew1jqTnKzhWTIlD2dtXt7sKXH7aBDWPpKRYc5kX/NE+MY82BRERE7TlS7a1va5Aip+0
RgDMXKPHWEbFb6WbUf4tkRbNYIkovcKCd5kEYDEW7GeWwtxoPU8PoGLRTzInAVOh737+uDazGoXM
M4wA9CamW3QCa9IlSllDu0Cm5yiHx031aRN8N3r1UWFgdlRP74n194JfccPiLjvFfJMsbOnyS9Kx
RDoqyAuPPTcK6N8E5TUEpZUhfncb47jHFBPAgAw/zel/LLKz8573OACJSW7LXARfRhBehvl4SX2a
pLoS4dlI8fST/Jrd8ATNcgsBrjnKJKw8pnT1juXnUB6Ks7ymsJI2mhXfLwCPJ4KX0gzQp8QiHiVQ
W+oss9kUaT6vlOFerHrtexhAmdlohp/7d8LCKSsTSwIA8hb6GFf7IjJ3Jt0GhZZpcFETRjUwSSH8
SpMPcwK2yFQ2/xoSWOuyEU2n+EtffaNs2vQK/43uwlYcKnUbvf3H1a7ueWfptDlMstQlUs+2Ni4J
GeRd3rB3msMdfJT7mhzkzzOMnGemDPsyaNmc1F90n0M5X1QxrT/26ACWt1M7hcifKIBF/jtZb72j
akJu0QCg3IcAdrWvJk4iog+sZvLjLFpDTxYyzhWRp7EI4tjcMVGIeszJNkWzWKnnSGuu4uJhvyK5
tGMniZyqVqkOHInvs/ugarhLCaUL5aWyC/bmpN/OiU2xBPoj2q2PDlJ0u4jFWVhTLq/2uXlmrbGx
19mvCE5dlDwjnIYdE1AJHZxPJ7W3wkUjYK1qvHP3MncsceYTEdmEyRvx3gkdGGfwRBhEvJupcT18
g5MgUWcYeLIiRQ0BMocNSM/941cNoTiY80S3xjBc6ch1a9GdyLNMZYEVgRLnHD/aHvrZ7iQoHU6u
tAeFfvTenm1hP/9QK3CV/jUCLM4nRvA4uhx32W6zjwOtjzaTJHoubXR4A/HCLYnLBeBGnjcVL9mP
7ahQJjJi9U1G+oklHI1uraajaHKdC6rOapvr9ngxWpl8m28Dx4z1gNvyE+Lt1OZRPKhwSMvCDGJp
a5X5uWHc3suz09SUD6h3PSg1OVHHxJkJinfWsViZ4dSoYHfgaD/wbey5gJ9UiKnTpliuXftqaG9V
HF8GBHGu5UU8uqmeNvfflBqV7vf71QbD5QrffIrKnEm6jqMf53OP4OCE164FSYjOfPA1rM+nVShc
bcoBgZVGhlaj6OSoHmKX3XVBoSiTWF8vcqUj1r/KPuUP4AIFQl9X5GN+E0FewT5LDlMz2veEtXr6
OL4yUBp9rYVwir8P1LPF26c6PxArINwvNyShCCEu1exPBCFps1Jqy1F6wsM6UKxr3ynBvFMbPSmh
ACdtQA3lXmXlE8jfD4+s94U/1FviktphqV1P2UWfW2DGCoNm5b+9dqF2qIaIstsxP4aD/AmCtnAX
jv6hTwsWk/rRE17pDsLw73IFu2mXF7g3rgK9T9oDmtfVceg71c7M3LIFTU1AXgt5oPDhpUbBeSIM
Zf6m6Y2Skgow5wFtG3O7vZrScicQbpwVjJ4bZDsmKFr2CsTBf+gYRlMWdqsjuOpPI0HsugDqVUY6
szlt86oGye+XD47EwIpF3npRJ6CE312XPLsO6KCm1UAxVF2vPSxklQ0jTZx9VkATphWrX2lv3Hhf
DEe3Xz98uWW8vhy6NfSDmL90zrLuspnvDuTkyaqyKjoFo8qzMCgWQR9X1PDb0RcPvZzYIHcgywVC
nl9TdAfx1x0O8TMtEa2BCEhLTnFf1lhMZGYBmEfE6HaLrMW9+D9sijNT7yNgHXO4kjQXsZsfznyH
/ieB7vH0Y6Wq6kABoiTG//m6QIG4O1ihV09lHzIx9xH6BBeFE5GRm/6Ocde37ynP1b8DQ9PtEsNT
v2tzqW+sXJFmHXpD/AneFwkupRo4lOnh0h5v/wm15XvTAbynmA9v+6UtIryYoau2mbignX9N9cFO
o0uTzq/MDY4hkv3a5WSfS6g6q8NxcaTHJeIozrOyqsvypvFXtx2+N3bUwQXOQpisTRla2NnVyH5+
4hb25X76EUUdk1wFbp5giQ/2Mma/V+Hw4lUA+gvRVRBw+3zLQMNv1+43DveRjcntRtSo8T2aSOVt
zfFMpp4Xdbqo6K3vc4N/3X7i/uAwhsJFn/mc3sPn2k3f0NO4HsEkyUAPnKLNv0YFLqpJoLwJOIe+
LeoJZ24NIJeJKUynh6bHXfFHYY4qylXx1qiIJNTQsDaBBvyD5FAYClm3FnwpbzelXjiiQIJMYPny
GLaQbWP81GUlsrnlz3yZ5779AFEwmtcEibVPRy9rP9U/YtHDWziQURb90XNWQj4PJa/3NyRhtMCq
DkMYHTru7Eg9lzKbMddX0jjA3oGUGfCYBUh2ATXLrf/TktV42HRxcHag22mAUN2SOFkVRsgiFvan
+odowjOOSIJXRRi+S0xFNwSEJiQMzSfbg+HbfjaCXDKfTK1JamqJc6qBHxTUN8FFPGSuJuZQC//t
C/UgWap9LyGuF1Zx9i5aXHNB7hFAf4suYuNJzVfZpHb6wmRGizPGVGKDoggFQKD5/xS8+1W9Hqge
2ZpNq9XHxzPj5QXti88LxZl+El218FZSCy/liQtN4/e4mao3P9uZ9x5nJorXJvPdaFzfnJWxKuZU
UeIbeAxHhdc3+NCdW4qTx14stvctlLfPJARZ40FagtI4WpE0/VxgjVlkdyHwSFWGv22PkOAu+aUA
b3NztuZNez2jk0GKqPP40o0YWoIk28Lf6gSuLMfadV5MabeO1B0MX7KG3r3ovCauMBUqOknN+lvA
0f/oy6OxNTudH0fpipbawN68C1OLSShLwc+zU1wcxDsn/0UEj8Z5b1yYSU0IBb3WDTxWRV833+XG
N7FEHkuCEgtZChPWZONYmLvQopvo455FhU+qkV7jX6HXpYYgaVQ75rdSmtR9CrqpBYgVLNGCcu4y
5OZCJ8dN9cmBI4sbLmCtogoiphbSwPUGAl9kEsjPG17bacjVBm8b8SoIsro7T088gbz1dwPiV4pF
V0u8OxaUxnT6y0wZcUIw4xEJwYA+itSE64oa5x0kiBQLPCY9IBrlgxatTDmCfW/mP0zE9Xd53IWf
w+9xNybzpc2fMcgeRLP4xdGxmqOFHf3SLDw/IuRvNl3dSfvYwU/S4sYo0HnIZSXmDpDrswZTG3aV
3yGTeCPPag5nzow3iv0JNzqJ67DqX6jlmfzDQN02uIYVtcyRXYyIyRgZhbAsocb1J/b/lBof6MSn
oVubg59qvSbRh33iYxiOr5jhGyGghL5Ie32hqvqDEnBwLWB2kRl+wWCpESWJWNxHi450ErGuy3Nk
ywc/pIaLsFiZ0YXuCdSgD/V+xQYGHX9y/VSsMjzmhvFo5NrFLuRXKGKYCuSiJX88YoYGqRoANIdO
0VpQdT5Npw2tVo3f09dAB2WmiMLh8Yun5rn7hHMjMrXSk9pXLNjg24cGsHlfEUFiQPY1vtKyLxFo
Qfc+2QFIkIKAsOPoXuZXSoJvPM2xtfy7IQn0wDK2yyE1GZTHwcqqnNQNTG69aN3q3SlauqMGCsSw
SvZj/mXWcp1F1Q1bxBaAiuaYG2RpW43ydTthbJR16/JGNnHP1RX7Jxm1WGqV0dv/YNKSagKnZVCK
e0oxleTNWl7PN79SeTqCM6ZWosQTF/7NhxxdvRWg1N25pXnOdpweZ0vVzKnRxtn0Yrf64poQ8P6M
tTAWwW0oU0Cx8zetOCupECH6w3ujlvXrcNxtA013kmxpkaTB1XfyYOCjffNUDQaK5bvehhK+EIye
8t4PJYcSCRS7HULKZPf/VjCn9gRTBN1d/MPLpBPrtgqFh6lfnGH6FtUOmZoDyzfLeuLR4T0XHHV1
T+auw7M1pcyWrOWzFvs6p+ihbHQTa36yZjLEpKdrmOClNS+YBtoV2LsETuZf9lQUzNiBfz1ISY/E
pTmsNfqFbN2/AG1RU9fl9VdSc9F7ZPthfWqcnLs8atv4rvFRvJMAPf0Yk8xGxjOLw4mdbXhgXLuU
zulYbNom4L+CeNqJPwHMMVtrYGu2cpN5pD2DyVb2XY0wbD0Xeqf+iz+4cfDVSTFR3RVVfkHutBI9
9xcZ9sMttx9TN7e9+q0ZwzyW2AjOekDyaPbrM4t6S9tQ26uxVipAA50lgPjR3sxzBazxvV38Q0Y5
0/fV3O1SHmAT1JjhRKd7IvVv4SMicRuuHXlukyE/5daCkSjFbzJDPwdJTETvywlPhwXV38r4iHgU
0GcoT19AxfnBGySNz84ykCVttVMirA4aYxgRlVKlACIsnxD8Lr3+Ixvn7TvYENIRtnKBAd1Y05YM
0fdm4Q9upi9HRzPaAfdoMc0ZRG7MU5Ma9pqDSsI8DVjh14B3KoNIZaeOUScNk1Dog+Ww5TRUFQHX
32Iysr3B1Tk13ZHAr2zuWpX6yGJFs0VMGgjHBFS3bjU1U9BwjNwTqcta0+sshFf1FDvvzr81H+SI
Jh4+5U8pvyU1oypVA5dzUVx1TgaFrC7A8AXMGEh3GNqoaF34Sr2P2+k8kwE6JoVbQrRqHOkZgHvB
eK9ZuPbnibD44cBB1EIN4yDe7vgr0WlFXApgcVukmttc/Z6C5aswSxo1UiI0aoPN+/pShevTRJCR
RPgiyYTWPBR30F0WX+SgFLgsN2f1AMy56y8Ys5F3L0E4FE3+xt00MhJjy9gJxUxwjLmWkbM8cytO
Dl/hkjQbsxF4CgJRYcJRujBLyhm4Y1dDDXlglmo/YkjQPlY1QuAZjpe2ryes4f5egqFldZH78MQ+
pt1XDF+IwEgSosmhnRLHgfo2dlPMoiNFnpY0hiBzvkzeJM5Iz5/XmR5rCm7v1z0tnlbZhksWMJvw
/zjP+nwip2t6LOtVIxHA14X5e37N3qJzi8WhY+7Vn5IKvw8hXx9Q0IfyvdIt9CxbtQ+gJGR+PVT3
6UxMIQKFy9ELMQ7HEbkn5z7hDqLyn1AzXgGOsaGPTTB/bRPjBbU9rztQ1Fd3xYspMkWsgCQw3c+G
0NDOiuh5F2OXFnCSPuB8IWng5w2+tTQFxpOl80Ccqh+QTOp+gSe4/oQ7MWiB4uMYRd2FqczWjtc9
iDejgl8OeyRbU1G9Ov6XDnrEltzKUHcctYbi1fF/tJZJbstiIWxPHQjTB08kqbgVrcxGZaPI4/EI
E7540CvM1qbZxFKI60Oz2yXZfTx488Xmqy80/O+Q7S1Ui8aiNscpV1crMgmDYA6sSlqeC8rJEmuQ
qZp0jJcSBv8Zj9NC6i3dqxuX7jW6knAcRrnL4GHmW6EQed6uRJG7U75LlpxRsWSHcYifVFU/iF/j
HH8aYyhGZ8k+feUHldv/lT58UzvhcIyipHZKXUZWfF4Gfa5QHRVLaWj8CfmN1fjXmlQQgMsb/+1J
wkELDODCmz3O45IAAimW/szm00anlI2fYpuQRQcmkxIGQ2Jd8Xyjm4kWIWBRMJMWPhWcYsBpdCHp
BEad14VDNvP55OEIbXEpot2NjD0ddR6PhrGoByM77CnsQnh07oAgEmcWM8abRNwfjV85GShLKPdv
poF3pSXJvj1W6rEFDeQbhjZ5zw60gbCp6Zjre4sAnWUGi4NPgb4zDj8ceDVe8yVsy95/LQxK0Skv
aBea2j5KQMIE9WpE30D3VvhSE5hxCcBQiJ7KyzO4tndmJbz7QKIYUlbwpLldDP2niyJBVtGzov3x
kdpajIQxr73kLNmOM/r0Rq9QNRn39dIGapCUtIAJCVDkIuxEI7phgkQFKmBpCWIa6ud/usJVsXFL
NPsMeVn7bNNMLSaL8Iqt62/DsYUf/6CWr0n+cyPgNd+fH2fMyIoYsfeFtxR9P9nl7fwcwnkFjFyw
g82/uidB8J2tj+Rao/6AsQSWN0fQiXM+/EgozJZd8GyzSweIk31LnMNsob4WOamY6emWlwwtskjl
iAB+uiwLmQozIIWdhBz3EVXscA9/zxtRoDLPbk3y1vsZ93H5KUXAeVqpaB1onWLkyyRFrIrcPznN
r5kDdonrMbO38ynDh1HDDi57Gg5aAB5HQzSTR2mGbEYegcGu5knQgjNz7oG4qGwoNsFfWsZXzqXS
U9NWMwg4BA1Gb/nK56xYqcyjAh039MQNTwQb9VZ/7kd8YF2S9N3Ut7O6X/yB1hT044cqQcz7Wofk
1dY7CCZXXtQa5bLqSfZaU7gVc7cVG95EQHzoIJpkGOG0AAWrvNuJb21gEKDEhmMJEBUBTVUJ9ZWG
GC3UaL7gVmJO4eR7dp5ldZ/isSs+9pgjZCP/9ZMrfoDJSZbav1/BIY9ctGlNFs6kD1b9gDnzAS29
aI+xqqRXA/QYj2wqnt6MneBLlu4yngnx6RWUGLzGjtx8wARhgVK1TUQIcTQHBUduhbvAvdVYNLOb
j/A2MViXfUCJGjfmL83RxBxCwOBB8VfDwlzBNUcyPEUpHQWS/29ZlZwstpY2RCKTDjGI8jbgo+XU
pgumnANUng2kr+EywLdUbrDx5/NWQOLQkRUu4NN5kXu64Cw7coQ5iLhStTKEOSnR7hIQwVRMPAh7
DWi3RXizT+dBVWN9OAvyJHRYxo5CiLZQUfwmJzywuRKlpUzDUAr5qaF32lBLSfdHMI+VaJakgIHa
5QV/tlKSIRV4AnaXzbHtAXtZ7SrUbBOYObKJH1CmQt5zi7B42H2322zKdmCx7QXK5RK6XNc7RNLx
r4EoTjSmZ72pcMfsen4825DOOpqNWdUpXHzOar0X4rOSzmKXbc6saHQ1Z/gkDpSOKFZK7C4J4Pn9
5rBuG+PeWdbjybXZp2TAR5L44XHDP7ZnkrZdm7KjpizgS8rR8OEtWUm2lAUGZcAEnXXh08UAkf5z
ge6xr7DXF2Wl+Hf8Ek8QajZTga2G7a4uzadc5Sz5jwZWweDzE4REA8L9gMzgGNHPue6Or7JXWbIp
grLzlvcIIE4rXv/8/7RIcMWR4Vss2aR7ehK5VrR5Q0l8rVJNLbV5keneeKUd8bPFL4X328YA+pRS
3xDitkt43Ihq4nKhgj2DeS13noxowEl32RPMqxbbUxU01DLWysFchIkc5bXw8RpJDHq/WlMx6iOd
T28yHdy1t2Z5xW4dIRmMxVLLmgOtljnBhNMa3iTu3phBfYoaQKgVYrGg36yl+NW3MiwK3VYB4Lne
62C0MxDv4nXwZQ7A7ipjUjKRSDnEThBH3qqH+0PCT4T3vqj2t8YJ/wouxgKP77T+lS8or4PSkHTx
3lA+qiuz0o7x3v34yhLjhlRbD2VhMs0aavMf3GGkQ2b8ip5+RnWad0fRJlgckb4z0IROjStSp5KM
mct8zG8IsBuNxfKtwhWfew14EZjB0oTrTl8VD9glpPqlosAOSIHPA8coDijuQMevW6KNweHBpWRQ
caTggYz93y1PFbnRY0rxnmCoAZtBqp5SSW9hwvVb6CJ8mdEjrwSd3dPoOdyXAVFdTboKVLbiO5/+
aZVZ2Tm1pZ2AYd46SPt1/g9n9R1WxoHAB/sUKnJWdIsCvhY+jpWbHN6WszlSkXbiTNmMMLteF3xG
3DmRvnqMXYjiDYgwTOS4gpK6dcWXAGaEtKk3hVAB2U6Eea6YcmrR5tDYt4tghxBQ5iCf9Ce8yLFo
e7Ez8zTXFf3db5SJT3O4IxH0PBKofMSYabcOTqfSeqFDgXKIhBpvt3kN5oOGUVbSX4T0Sfd1SnGx
zGG5hDwQSHrjlF8Wq26kFzsBn4GFx0RsltWQPXDr0WbtIny/uB0C7c3cCk246jw7rqPVGJcTK/Py
k51fIQeId2Xc2jTmDyayK9pkP1xapX0d9IEheqvBvgO4EzqbxgqLwATEL91DT2jAaqQE5nMsf4su
5RsHDzwGNBBzv9wGEQN+h3zDAX88MKK2yQORp3ar4F/rwLrsA7jXJgV3OTxYu/Wy2Rha3ijLEx8N
wYVhG4BckowYmu7pD4YbAfyz9F31epnw7ClhggSCSHJlr2k8chRLKE0fO0T/fE2E/yG4+6Dbegbc
VagwLmIjyQV9mcS2CA==
`protect end_protected
