-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Mez040IzryVDcQGEY5ve1gcw937YNlZXUsPkA1vdqjVOpSEG96d0ScA/7zPXdDkPJbmLnULP7Yv3
vP3/yF7t4oWkPdREXD7/3f3l4/FGnDaZE/Yd94U8l69JRMqm5aO1ZIHY4OJ5KknySMubCu8u6Dvd
iE95Hc6Ig8gP7jJufWFE9GrUGXi5wFUTvWH3APD6gX2L7YpWtz1BbgP7DBOEfZxvxLvg0rokcbRc
z1syRZn9tWkWxddA9vT1GpLZga/E5AnaEgIV+V936dsZ2s+nJQuJQ9GJ01slL3NxYPlJqM+ciMXC
IcyOgs9rQvzYqFG6hD3yIMLMS2lO735NjbKKCw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 45120)
`protect data_block
jEQLNx8HQeAiHD32mNOXkrIbbv1AXaMah5F5SunqwSWrafZz+zXgmgOWdLnSl+kdCUS4tbOoEs6i
lOrO7Mb+CDewOn+nTdMbGs9V6/N9n0DCwGtj4ZLjlN7YTVj0ays7AxSQrYUdBqlzGLHRdyTdzSHc
WXBmRLPmhoVNWICqEXJHzfQENgrEZ9FX/EMoPnZUQan3kw5ADthfQonpATQZ5uerfv1NIzuj1dvY
A4S8FJ1XZbSoptIzzay9MZA0G9mnVP8tA6djanEQ7o0Tr12MlR+yo0lTycA66gD8ivPkKXnkKC1w
G5i/OvyV7QNFKR9H/ZtmiWnIX3gEkYwTA/WSITP0PDmAcPYTY/zqNauCcWiHfGJumSZoO8hKDoeG
UUBwxgh1d8RxksFb/ISYodi2Ui9O8tWngoal+BocMxXcM7JpB+NXWUC3EBmIoxCENsbsG31ZnnB1
7nS0eHPdI+n7ikXVw9QVOsMmaA3hUDPABf3ex4qxs02O/6wXHO5Li2HiWspFCDvO/htR6P+TZNXk
BwI470GTMXAs3jHrVfiF6IlQkvGmjvydqUoqYgxb8606QfiI7fumRZjDIeQJO7VIsyf+vkXtP8h6
0NPjfL00yy7cAl4vkOvD5hAqVLtYLKVeiiC/bBSWzwNZgdfSTkh2eV4BHA2joXYJwmmhCdZMfn/4
f+4wcVKdUxEJLw/DKqzIrcgyh7hjpGVXU2tBNTmuahHc/kQ61MJPHNsI5POe2p2TGRZlBRFokILZ
TWSXezAkGB8rZYkPJFQXCbPEwlY6wkdlUTIYUAxfmNGuI0omR+0QLVeLQvp6alOHiMICe5NI/r0p
uXTNZ5En8KC660PX4btPqj1RYLB799H0wUnbPNxHPz3GOqBZR3khThcvEtpUjJZLVvYM0KUTV+4N
3rNDWVMsV+6VLgE5092ssSxD/gRapD0P3e45kkhxV1cR2pZ6iiu0KUBZxvBxBU+U6osqVtrUmlF4
qIxLzex6hVz2o36uT0cuIK/Q+x0JmxS33fa/h26Y8PH2wwEvxbaEX0PTwuOPlw54Sa0x/l++sJ1e
mJSvcUtHM2YPtKboZOPcSqAxnLuOu8h5NydF3QjwqMOhA9vptnaOSrZtRzS2Rn2Dly+Qrl1GE427
kz6+sxkYTpBr7F537oIUBplvO7KhhEHVHTqDltL9XBqr6TNn0s4vvakG2sX7jwAcL7oF1ef6jZ2Z
GhoaMXuDdlj8d+JknWTwmrkZHbAQgcy263YovrBgVKXR+Vs1xzPCeY75hEy+yQg4T+Ep2rFmEwKS
KiWJE7lDxOtggngWlu/ZLYUE1JsaMTX8uaoEJqkbNhtVhBABJeXSGFGx3rwZ1pDYg5SQEYvA3j/m
2JVXVR5DHcStFntPROAIJCU0Fw6x0hFYXPudFwfL+V8I0OA75S0/C9yfwO5QS6L4XtB86ihKQPTP
GKnNATV8q3oVL+IngjRkUoDnj/3qP9+UWxExIU2JnPRGcY8GHVs/dy9cVFsc+1d9+hihaNkWjxqh
sDoAvL9sg7HSgUV19hR9PsoAXxjggF7wgEU2caRyFeQBUt1msU3A7vlh7IvHzdFRV1l4gWiFishg
eueh3wHhvi/Fd7q5cUK3SI8/i0ZlH1R5qduOs2UGhZiiwXhYxNh3j1Ql5LCh20uYAH+Ec5zLjl/K
7IUPqwmfImD765vpM5K8uaBofl/KnYA0YLnpL8+vZiQ+Es4YoC1PdwHnnUhtoys40ZFxxBvEGblr
YWaSrnRNZv7PGi83o67nXmDUN0xGmB0AOHuM1FrkGBgOEdZrDIAIYv4U83YU7bYqNLA/2FkbUkAB
0WaY5uNQtw3+oRt0T6fWycq4rnWQztaVFGX2HH6104ofVBceLhQ6L2PjdRUJ/LgsTWXKwbdNfBAo
rfdyo7o/HEJ2jAuZtbiAHQ2FWvArEUNN6+mR/chUGwhe8SKhWFwC9cKw+PEJLSJhEDMwje82HKly
8KBnbZ7U4ZiWxZJVB0nORY9nd3wK9aaXOF9/kayxiTMZIMQr9ecZk8ZksAEM5G7EVTlvR+Ki+p9W
7F5Zbr64fQa/j2VGbLPgFpd7daBq7SBIADrVcTTIIxzHA0WZtUldwcNllVKSB1Z/ZYn1YQQvISty
h4g3gyO+STKaDBmSr+SDNyEYe3u8hYNXudoteY0Iw7Gryu+REHn0Le6yhlXrmN4FJo1Knng5Qy/j
Ks0XZ/0fz8kBq83u3pe9cWJ+wgob4UGkbCPRnXbmFsRC5sYyjaYuaBhok0RdLNFN1h7V1BelI+8Y
uEVDMzHwocXKnPK8vTYopk6Bsj8ilG7K/sBTm/KJTIzFQOeaAmm5i7coMEJv9gBSbFMx6KnNnwEq
5JVppBOh95xLrE/7Jd7qfRvsHEZ9oi8eugMIdCzrK/GQuVNB6iUrptKwhKMA1rpcEUmqOz3r9YZj
ikn2c9T8I44RA8ZIWTaqDFPEiXCgnAQhgsu5OOrHDw0cb0xJfQXBFBKvPLwmsNJ5P3+7h2Vdic7T
2Oco0dboxqz8J1/5esYS8ZEu0okHRYU4yBuDsaV/OUVqtXXRkjq2o1uN92fQRgbi7LdgaSqQyctq
Xy9NxdZlpGReHtp7R23AIS//1OwiJ3Th5701N9pgjnWUAeUrgKHqxKCulqnj5JYTFzusJ4s3TJe1
Y8MbJmElfLAY9mvgpSL+PY8kJqL9mUm4B7ovgmiQLEv0ggQdnqk3XVZgDlUZU2ksDp/CzUhD3R9w
/9602ti7+MvCiZ1wO1hsS0rDRvuesfddlmd22fFj7uOYYDLEh5h7zSkADF9Dbygeni8AHPow5jmZ
IGX6zF61Gfuopl0RN/T9SmnHmpr2ZNq2nWFIztGhWZstvfamUfhmS6qvbTd/tTYgckKLz/saoL1d
OtvUlsyYRMOxBmWQWfOwcFaIi74xmcYjPCzdi7poYgK4+CEu9h9ru4RHUK0n7RncG8xcAD13d0hL
pyAz/FVYuz/0AS6aF3yuLAejGP7c6uX3e5rzZVuxBfMwmUCu79FuMhoAORpj+AxsY1HH/Rka92NR
zXJ3Jz8PEmIcNIlfZY5Q2qlN4enX0ScaU8rzYkP9KlC7atpI5P0tBh6TCWm2GjFrWRYlIHy8eSCi
wQ6XYc6HetMG/w6HFdqx237tjxh3h7+bsovpblfylNTAeCXBfRby9Nq8qiL+yOzqpFn/oGJB9EBv
0pNFjp7K5geyluWJb7wD2oC7Y7v5s+8VyqkUMMKtPMew1cEW7VvdCXSEkiVrrAwxJ0USZK5vFvmt
8QC3JKD4gvAB8X4z4b8kEcPm1n/r9UlATlHxLvCwIGQNFCAZGevu8Zqzxvu8oh2fSg72JgxYigSq
6ZNmYHzPvj/4dFZOgQiGSGvlE8kEBNYPMVirLo5nam0noSXgf/K12wanTfupTxrKnq49zFV2Xctk
BaQXDGHSegCZFiFE8N7mEdxBi9yabyuwXN/Hx4hY9rAyk4ffkUO1J+ebZIi+pDP0EALuv4QTrCMB
FX+c8L/Z+Be7kHm4pUCugedZyfESP+czWsZ/UAC+HrgOJ92GhlzsaHG8P3Z7GzHNWHc7VsM1AJAx
TX34pSyZz+SSY4JOhdQNf7OOUqEfPZ+TS39GlmoecDqEoaF8RSH7YiVBedAhk9MgdIqJIlCJ01oD
wlnMGgBnUjTaVznmjGRISe2Awz3EqS8VO5E5iSmnchj57TYzHHmG13q+2lQ5zkEStPyayacZz0mh
hX/XpyMU3VIT7Uhs6fhzfjtYfUoNc34/Fo+MdunOLXCLKQE6yW/Bpsq48oNPrhT+NOpmGtXiTiC/
cNvywGSoYNpd5zCzjGV62kVm6GfO59ceFjrmpHLXr3VoL+6MvKI9DtOpna9jVPC2ZdtrBej8Ig1V
K1gzx0xdF1tUZxf5ioppHcYGVFNcpqJAUOzsyv17gZN4dr5fw3SOQKtTT5p5EQINqExMmlRWjHlR
tmw+hVwsybDTjnaGRc6r28u/TkfslLcVLZ0sI/pESf/fPEXECSHgnLtFqXREbHqRXCkZzNVoATZQ
cgvxB3saZdr27PpGCiXWoueW7n3iNERDzFeMRDVVmaif2MjXUFxgBhlyChGl7LaiBfeRrZkNkSVH
P9jdwgjOaR6uOlYtarIDgv+bUp1psfRUKWcpYo87YDgWsuz4kDiwM5XZcc/+cAlEFEj9OCoY92zS
bNLHFcUU+wR3DzKPEvmSoOTCVJ8dc/ZLu1bGafmjgY5NqIkXutHaunCGMeaqSUJpQn7SbNsx1sE/
U667t0lPEss2QhOnMu5s+WxyPpMwEKqCOM0A4hmLNe2pom6k3ga37gsA0s99N9ZqxAOWdv64pxRz
a+oGH0G9mWP39w9L05HuKDtW6/eIGQhPk/AGZanIyAtZ0G7szcwws3A1B47y1p95skRqBgbdMW3I
iPBCk6w48dYF+WZ+bULDnadTk/7ZoQEcu/UAAWlVDuxtm9k6ueNY2heGR2Yx5yfFEMB7/bqgbGe2
QIuVol3oWUe3t72P7Y+U8AgcbQyQe9GYvvmT4pcE/ISagZKDWdxmTaO8WubIvsLAD9Bt7wJyxDCh
AsMNtZfhbnR+42KdJkf3jD/hDUC3B0iBJaYsDK8z70ERjI8L/zoVpHNAUwx9ZL2usB3KmoR5YTVX
9xxSQlGbDblvxwuquLi74iuQ/zVHmt6tRwcTHIWDe3TrFVVFUQ58nYnA5PY94+ViEOz5kXAQxyeI
U2+E6OAs8goYaJYG/y2EGoSE6AV6Vy99uvufXWBu0LY7t32Kr9lJ9TbX/HAkf9NyCsNXzS7GqpPV
TBDbDwTG91EsnRalgU0zdJdyZK5Pc/2PB0gJWnyYAIjJERc4G6ienI2Qgze+G53MAwwV3HcrLHx9
7wRxHOapAKZKDYkvzCBvaH4xSGBMbCSR7PS+JlimIY5HC/+nW7uoOe74HzJgVuqmalaRKL2Vr2Hg
JfFI0NV7PUuEta9xnprr4dv0oMCqH4O3Im8M3iPpgySHmQOsqCl8mePrg1ObPPaFXnn5ypS9FB/6
+WdFNLCmK1OEeL54zPoRc2GJmL0Sk9niHvT0vhdvaQAYsjrJuA06yH6MoTQPOKSrD5d5sOUPxS1G
lXNnVxhcHh/iZQFr87LWGunEWFjHXcBtk6qaExhVs5wgmj3k9NKq7Ney2ko2F9tnmZIDWQPxZnwW
EBQQTvVYNDWVS5t+xPnBR9ic38O16Nq4mqxE8DKGQM84Ak6FXptXcRtsaYLH5+MrDIkuZspE7E5t
WWBhtG2KeUSKLbNqWyPBWvbxKQouyg5EnT40brmv5yd3487UaXLXaJI9+IHqpRQFDMaTqT0fLqf9
CeIa15I1JwIqlP2FQJiUp/JkuNNVjSe+aj1JzTcySe6r88MmbC9e//dMGDN0WkR8RT8Pa8atSiZ7
S7AMh2vwkh623fFOg3wE058/k7QRnR+hA1o2avNH1Yg/wWeNvcLgEXEgv3d7O6ReeONNauLSt0P1
Xmu++dsJPEH8DllzHg08SvPEmj/NX46aCMWQkTWUyBPWRGqg2M5f7P1rM2eTtF0N3p7fqXDIDmOY
p9QOU/3ySI9koY2hX6EAaB4APaiAko3bKbDJMaArBAbxKeH9hLqU/kES9GiVPaVklZWSlay03wy0
pXo5rjUWktR0NEQNwIJl2X7BZrC+6vjhq2tdbKEY5HZc+o94q186eC7jbC0EB63yPlWbgd04G18x
aJBXLq64ptEfnyqmiwBb3diQxW1GqINXtfuYaTZa0X50wrpjeZgctde+8ali6h+0V4GwYq7DvLPp
K+rTYk8YyFYCZNV/nxFyPLNPme717RJtQntRVBpJqaPnwWn3tXBIdmp5+ZQHTcqufvVBm7oIt+mY
Az/NXxv7re5sTxy21gm5fUvMYTSBskCskgZdpyRwTSJ8/YmFvO40PyT/r718hZKT5RnzsUkM3lNy
7LY29g+NNrTEmsUbQWopAo7/SeGBMGy4eF8TplPKZIsDhRsoVPNhuzZX9dh8PxfcV3PNhnCGIiRc
/bbkFPRsBZLD0Z9FAKEvgrb2MyOZjJcFM24Gi1d5xmBvZ7hUhiNKF5vZkihwf29Zh6lJDbOA4Qpl
HGWAfi2Nw9kEvxoMg6aolK+BsxsQa7aivdriwPBaChpUE/jFwfR75EAhztvuWZcwk7NxfxoLtY0h
CVjYqdI+RybGTDWo8lCQfalpcgQy0YYctFE9JLg/UwGrcol5AY0qyMdS0ZJFm+1GMGuLf5nvoaGv
C7MkANmeVySrizfBrdwuxS8zKqU9U3UtXlCHyqcpHuP0TyFnV4klAjeTfIpsF6/jURFDWT9tZbcx
mh8tWp0Bob7rVv9L/lXsVjgUihdNW+MwQ0pzzFsCM5TWG8RMhkhpp413ajBrN15KrMOdsoILd0ne
GOFTlj3peb+I8gaxN6piENGu67etOPfv4DopmQ5l9f7MXJQiVdjKascqPwIUbpQC+y/lRjw7Ckaz
lurKL0pI6E4x+sCn0wsOcmXrx6wTolSohdPFqUHkS2h0KCYEI80oitzjydlTDbR4J1qO6MihE9tK
VW1l2CE6wR6FtQ0onvz3L8uW4KdV/2NNNBSACXEIxQADj7ejOcm0l3+NXHkmL3CXKXh97WkOftY2
lBFqPMwTUKICPwXSLtNfeTxBmjoNW7PB0OUiAhjJomKoltI0sp20HbuEJ8PBGjEShi12d8JEdTIu
H6MHY0mur1ESW1Mu+ZKfRusaYT9mY4mLVHeJ8xEEClDTTtXcDlYqqlPqwujRS0jUfuVrSePVXreR
fCeXDNUVzuo7yZ20bUoAI2s66wiEJXCm7YIaeDtDAz1hvNo74F+O/T+jqWlF0FfcF8nIxeZ7Hb46
kMiwOQ1LqAtLnaOhmhleFRpfgkE3c4WJqB26qRaM0NKc8jtKODaFkQyyJktZ5ZaAfLxij99YEm5s
XfCI9rrueSPOEHR2t4CaHFz/9IVQ17QaWI9NNqj/EjnilVAyjqu/dRf0WBGHI8/kn+r6ASmv17RV
J3JLhQce7mjrm7ZNnRWAGgtZ9Q1Q6ZQJDDSGOC0uQ0TFqQN3GTIiefsQjB55QBmGKRwycsSwtSOM
m88yXutzhopKcq3JHBXKv9Du4GhE27H1zt4fcJSEufr3C+ksMPkz/T2KeeI7hNDdRHHazChrU7Xe
qgr4HNCmdrnpZf9Wig9CQQrWaSKOSvNN1rC/nedX1fKz9qOYOe+zhaoyVTMY3CShnJrXCPUu1z+M
Kq97m8H4n/5wPIrA3wQE86At8Cheih+h0gT9Cjwi5RBL5+yJAFQB8Xm1i0LQvE4AZUYis7CsfjIH
4VmXaD96CKQqtVutrxP6TV9mSbPZ/QH8DT0VlC1pEPQWbXIR8z55/QBXS8GVdN9z+XJMxm5dR0/f
U7FpdFAaRhb7Sd5avsF2gnhnneEQ+R5gOIi/FZ8BUjaO6IoMDHZdj6uCHo3SUJfhpsfrzMrv5VER
FaASUieC8YWYnSXNNlGOr0chj4GirfOKfLYuRKr5P5iAw8IkXYvSDqj0x/jF12OknOzK5ql0+Hrv
XE++VWlIcdk+1hiVJ9QrAU7R13k6gwwAz2kTaZOhBZw1dqCh6eFfuucGZp2/Kf9rsc5DjSBMf0lr
n4GpBr4EHh0M8nqjvi8dNO8+iN+x05Uu16rEGKuTI6asMnk3xMKwuyLrOEawZZASdXqlIEbtSoEo
D9upfKB9D/OaJw+RCiakeGgmBrPXRX1/0iOnM1HfbpHyx8GCyzeY79PONri34SoTVXaNDAYzsh48
d2kuYzOaXWPiInsoMNvt0L8tcSnvE/cprU1Ta2XZSMClgiqBra6RsNWEKorTsg3V/5WO3pq2DAKQ
sm1K1+z3DoZu23XPu+FqxckZbEY8+4++52FL0PGN4rx5OZ6NeJgMQArV/iDv+J5mlNRWeCGBDbMs
XDX99M9WBizbx9cOS1jxlM400D9krVtlxZ3bHMjQjPPvxJWxZPyMAdG2Fx6eNVdSJRvJ+Ad4VrZ1
KpHq04N/oIBnqpnJW0eemERoKzqSeEGyuefqzcEgU3bRulUYIgRmS44H72EKJ2JvNZRa9TDlkcVJ
WyTorVmZJQ6VcIXfClf3YoF8igXCmwwLdZnL6zU5AY0AHmBb2+sRYUqeeIEcM4HcAoxhFjU9Iq3W
KvDc/KnymfEhyZ966yR+keTwcNlDis1jF+HL4iqAfAJIHg/cshQvB/UOIEHZxCEt7zoSJkfBu2H9
jV16n5h1fQaNYeWC2mLIgAs/XbHkpVDUUxvjGT1iLyex3u40GM1ZbMBcJobUd095j39fQ1PLjavo
QrqsgCb+nUJRksY2LLd7zVVl0qmLoB9BwI5jthmw0+hKfPt+LbhMXmwjNRLcQKWCGBBjjVkAsjwk
HJP1l0P2xvm4by0Hd9eDzJ173wKo1vSd0+M3CtHYDS//P7SWdrNpfbQPqXVA8oGdlB/R0s9J43MZ
JqF9KYc0ZihECxh5bxbJ4bM8xdJmvDdg7au85oePaZ5BPFJ5rmaS2dY2EpUejusk0qzQuoVrxzM2
SXWnduc8qyF/SkYzMgbckB3lsveokIzm4GkSPLbUPFq4MmiwJdymOsQe0dhJZ62597FhjpiFYOMp
XBijJ8vpolkncAArnYt2LGSWRuWZNS6qOwb7xwwNqwXy/SV0CwagTkABiAKUq+l9BtcK28grn7Gk
AFNP8T8ApSM3/DFayCQLJWV00n/h3pljyHrr542NBzmSdHLawxKikLXxOxRknfNv04uEvUKnsl4B
IA2OozR6vR18hWvR1DF3aFgSISsd5A/sOBJBQbltNpkqh/pIOGGdLNnQ4iKhTtVx3FIMEPBXP/XK
zCCo9FBwdONyfYgkxl2kA4ukZCbr55LepHkaL5r3qJpRuYef0D51t3HZ3yxodC6uOPTrlDG2y3CG
UMGr21NgT8aBkLDni2sclIDKgHkZsTmTuAUtZEx+KnsyU+tD4T+XeEXT2X2/tYXflBSvcCHaARMa
yAE8uCf9Ec62dNjoAj3fD3B/2PELeFta3hNH+3qDYFFEQq8f0PkdWvn1RB+1nJGpMWrUDvOEfY6b
TVgWyjVpoxnS72V6hT/ZFW0LAIVygA8NqefTBZ5nRvX+Ue+Qq33RhUMdSmgE5y9iTux3D09RGLDp
KvLMW6Ac9Q7DBrncRCOrJSbw+zgO+MmWi/oaHoVbDIKe/lLCb0jjmxMtti5PfW5+0RbbhQdwSrme
X1GlSFI8GmTHyC2yNNKw97Hs7aMxOJbO7vuhFdC3FncniChBymHuKqxVDqFDRgYGoidytNMeetlo
5Mp/HyEFhAUzVM9R21XwKktR7ReNlKd1l4L3NAymlJ1jT1Kne0Gd1MIBFTKoaHHgbhKKk44hSabt
GyttYg5ltrob1dmecw7SrNTEz1/Kw4Bu3AkFA+6HpEJU5q3oE7Tm58QfMfunEzGBtAdjuZXoz4bO
uuDispUf8haA+PNSBB1Ypx7pzEFtJry5XuAg+E3cuOBOpyEuD0oYT+3Qyesy/QrxlF8FFrr+WN/I
MlXujNNh0K/FedeOrh5lJQ/Toae9wcQW/CRDW/z1V1XjoT1MRLAM2M6XHDnqq9n8J3cd1QOH+95P
vvR5tn+PSrKub34Ak9ilbP7jPPwWeLGePK6sYVYJX2uvB797q0RXnRt5gT0ofOOcQPtTTv6F/pYq
BzCgL48IKTjiXXfC89+Spg9kcqrZqtckGZWgOIz9LvkH9Vml6t6Va7nl2dv5fYdi9lZmkr1Wg1xE
6/DEZ3KXslVHBIt0Ea/ZEe1nzBCmJA+YS64hrhkREPgPFeMHi33vGl+fx+STqvJa+4xOngrfXSeR
zJWdZKzZgx+6o6P+31F3R//hYUEIFYfLvyZzkH5M29Wfe6wvRqLw1sObqs5+/KYXY80htXsR77Us
+x55aULSEd6fA3sIrI0+v7Y1bGqdyREKoLga382pwMHwdDSpuVmDs9fHLMGdk75Qe2Bd6XjbqiAU
1ejr+IwYkOZDKj6LzpJNZoGlSTIY+WHoCyurOAO0ZEpP4ZrdbhhHVXra8yk+4OiuYzzMzo20eZE6
Smf6+iMkQXEWFvnQDFGvPFNIEtAG0XCitFqdWYQbAldncwHhjFl9F/z8dSAq6A46skK+Zu6YGTEQ
iHp7BI+9R52k2X7MaoA723zDEBWnJSXMjv/GeKMcWKV/XYpfzs/hT7Vw6zjZu/U/1UeSAHErJEc7
p4vHhrrwP5vKrACaYj+Cyvx3kFFCScZ8F3mcCIol0QoatC8/ZCYk2Q28y+hmf/XneAJyZL0dA7X/
VoNnt+TjNSl+/owazEZMLTeBY6UVB+C6vcJQqXgIRHqYpaM5Flak7U5crNa2qvNnHY+kyvuuf+Gp
Uzxw34YdU2nLv/D/xX/O7z3cVp7UDIE7K5lHE7tzsoAQcnYJRib9cqPZT+jHZLF7Sp9nXjl+VFCD
HH1bLrGIacuMDNFbVrlNVYOnpnT6JaD1kyPfAhM5cP4W+DiJZ2iusWD05fyeNjsQZ+0Lag72prDu
qMfElJRNg2RLLiHbyi2xWS9Rq4nP3l02RImWF0fvOx0bLM8xvRLkd37v580zna0M1tyOAYVYifBB
kC1AKJWfgwtBz+d/rIZQw+M8N2IrNR91PtrKwISftPt18H76YciVzrgz31+OMR6lQbeNbKZPZh8Y
beuN3QZ+fM/QczK/8Dg1SJEXd837OWgzy9XzFBI3FYUH3SZZifbqPGYdXonsNE4QPFCeaNrPTOF8
QwReePoPGaUbVhrgZI4Hpp3t80ekB3DXykdHSsMmB3k39fReBIkUTO7mXOEQPGtKL8bXlVJh2lyr
kTkTK0hfNZB/0BahcBS62XaV5jtXGFRMLOUCBjHnkbBjkqYZJ1DdDDi+R9nHrMRp3iVdEvld47DM
RHpTYGqae6TXvy70K/S1SrqwkCq0WNfmr0kM5FJcsTZejxakGsOcbDGWTWJ3dyWTj731eStiyM7D
bEv2eMBz4pP5HQ3Z0H5SZo/QAmMSNIkMn07koKO2Tv2jqjCNm2rEoa7EjhD5wnRBhz2klZ/l///F
NNVyuUanP5GrAZyO8+BLcqDDgKdhrGB8Ex+rxFJbDcXaaOucJNnPxPEiBFgQ6lCkd0YkXhrR2vof
V+BdcgrqFl0WdOchZKNmjxDneCzCiZxAU9s8SOKrsE0DvxngCXtr8xycBsFkJeIhRPVOhdXG2AgP
7YOP2hkc+bYG4uxHiPVYGjBjNwCQ7bCzWNGpBCCxdlL4yof9jlhZknCXz1eX8niBmmqnc0dQDX+e
yhKr0lRga2zFm2/oTY1Ox1T+t473664dcy6SJ3a6jB/rfizyk3ybNvRFH9xg/eitOhLkhfac9d9y
BmM2zzNtbziKdFdKZdmrrJSSAM6kEEGE8Jv38eW1Uqo4MJGtcTdMJzGGMlUwsTsuVkQja4chRXR0
JZWWKTLs3mRDYLBPhlPqsEp17OFubOLERqmThXYkWuWPQcoXjKVjD1QhABOsGhGxd7Dc53np0MO7
43LvaYXAS9oRrTwQPZ6uJ3uPhk9oV5kr5zmsGpA8egwQanWnle8DinM6uJr2TlnHrHGeoCx4RMrc
c5E2ro7p1bVMktQY/QvfwhH4Mkb4x+HsvJI0UpASiQdN//j3ILsBOm2vjbfBQ/zxbadR1Kr8Vxrx
HZd6bTRm47MrDR7EqSilopYYM3Zsa028fozlbG+3vnJUoWp0rlaeSJOtsUF+9xQUHTL/0yIlLprh
HaK1vEO8wdnYbecfkE3kyPSrUT7kB8TwpIkjG/Y1HaGnxWa2GK5F9kVKax6cR0uiXoblCWiLFDbS
PsdTvllhrha4+nVSVwbEifA9B6b4qYxvVNg7ikBh9cEsiqTjKyfCBXNIRJMftrZXO2fXZswPgLGl
MhGTyt/hzCMYp9Sk3m9HEGiQxfHGKgHzR1AX+xuJh+vDo4p1LJszERIcgaYxgJcZNnziTTwGsord
iq6z0hygq8z6uEYUwbpvOPKn3th5QyVye0HV1r/owF4Ap/1fpRADKU6BoIDzZ35YgmNsJq1iNfYW
tAAg876Jk4SzBKZX7W75KUMJ0jl01PPIP72s3LFlImoYseq2J+UvTR/LxD8RUJ0Tn5AaeGhZdFhT
SiydLSko/vF9yq2gpkrrliDB+w5vtf3AgXaKzqJk6HE0fG2RbHvnFY7Gqi9s4iiAaZlQ5KFaZvMc
HOWB14w3GpSOb8lqIDtjdSl9ew2ISWhqnKRBgAf22RRdMIzzAJf+z5i0iWDNRJ83NZaxJustJy+A
El+2wvUDcQNZ/W+W3u/eDCY/FVVA112NtbqAr7U95ZQfTsnueTX9OZzyUx2LxfAGrE8HtUKvnsbZ
nxz9uIshvgtYLG7NQJfGItF//COkMKSlkK0YD7KlKNs/5SxfMPGUGr06cTmgNhclRBLneQ+eygu0
srztkG6UPfRTqcBp/2kP/Dg4NjvGnUkOXKe05bY790LiwS6aHTMIkGZPVOTjpQxO3HUa28X96NJV
2NP7ssNpFHAb+EfPQcqXAX6S3Rf2V4qLH8M+6TzjTUXPrybnE3X1JfKd5bdZaNq+RVaRXYeT6Hae
TOzdSrcPH6AMeqVKKyH6mWpfG8XyhbJE2W10SyOUlItJlps22Tj+bVRjGW7/ViPmiQTwVjh7Ik+m
fZMFIyVnk0ZZidzyYd3t8bbHQmqQDz+IwgxVVvXktAhGezsBMaoaPdWKgVVeoSa1fOlCdmnoZxFD
Ya6zzVEbpaGCqHG/MMo05GabLl8CxgWujWQLQv+eaaF/ZEvEhrz2dFepx3IKaP/EnA3TDPwpBamJ
lsUy0lTQm2wJxC0ea56Y0Yf/Tuq/p0Qut3tl43QSVI/aZTMkEwzTrYWGhqxYSJ+QRjXR0HLGzH/7
sCqPRoAL6T3YLsX8aNIZ4NUVF82P9jEzpGfI5941A7QjrmDBWO+2ILl/vpW6TOKQ/R8rtnX/PwJs
gpJxbTBGTfB51FBoxowFJBmV2FsuiwjQCTqQPsWKFI7JS3V+O3zmxB5UcAY2daR5BqLldxHJwCJs
E1mwUCvBqFIOf8MmI48WZeWbwfmxq7K8LnVrJWogap5oh4lXSTVand0+q0ezETiJ0aQINXxpeA1S
wp8Hj9c9phkycug9T4PIw6nL43YdWDl7iGz70yLTmAJpwVnF2pBoX5f+BT5jTiozuyEtgfH5KG/w
8S+yJgS92y0lOcPqjs4trKKipZ/9NqB7qxRlJf10XeRv5Tqgu1w4vU0//SWQsUKU3qCTGxdp513W
YaU+BfGnQ9M9ryR9E9x0vsW5PxABKyRi6RyiMdSn9a2vLsfa7TuP2bFsanKpjlYLNCWEGk1qxkbi
obN8CJZgZ4T9TmOefjF10CZaS3DguauNRrFhCpU3LjQSkRiYvcjnvebm+40rHY3UiCOXfdN/Q3Qv
cJ2pQ3IeIHfuOMyRvAzxp/CJmgbwd3X714pL6jyCQHCpNFDheBMldq7mHJ655oAZsTVjQyqiwEKM
9B10WxVB+BRwxlgIAKsPfCor5e+esRfQCy4rFLgdjh2oNo4jV0nv+3rxjyXxckXcpkDKXYOEsMzw
mCjMKgvVb/Bk/UY1s3ZbhcEN3avSsWvnpeonwQb+op23LG/7QIIC42czrKcEo9jDvlpobPrRAXHm
gHuC5cA1AJ2cOTngLOq/8YD6+8JqczMfU8qHjjTgbZ3gm9CdFZm3EK+rTcD6BtMdR8rtr7NDvVQ1
hFewMas2Vtu5O+pKBHit/2lUMxqKzKpcdnJU7/8bwswagXI91/YUcmOa8FQfcWnCHVWlQtdVVRGD
Z5EKRG4z7a2JNFZB5AEl+yCAKlqhrJLFdZaWoJYeUY6r/2Wj+ECbBOK5uNBZ+h44Wiz6B5p8IpxT
X/tq9vD1vnONpmbuZ9qpru0hFaZ/DLJ5RmS0/6oPS6t8pXlD79fb9J+ieuFP4THoBR8NoIY3mcVW
ae6bhu/l2OS3cYNQs6DEia6/zw91QFXoKUnEWtE1thb3Q74H2Vr4BqxMK8E+G51DBY71Hluy+BFs
IRufOFw1KzOFLZzncZe0ZrH/+Txe8x9J5uNy3yEhtBYHZrz6GOb95+mW+6DIhiN48K1GSVH+LQjr
yr45C0FFH0cybJ8l3Lf3KHpVDcV4filDuArL6bKqYoOysowSKCuPd21DZfd0+ru5LyIktKRvRF+F
f/gN5/pZlt+krqt0g0RsQU+6FIsiWFUwZ8cKB01uuJaPjicaPS1c1GceWbCWpgEJrhmFn+lxNIEb
jjYjFs1IEmMiXSAwlxxfErxLA6p8P1JI5QWB3BDJLs2NkYPF8pfRSa0XYwI8/C+9fDLHD35VH/0P
7BZSmUw0+bFjWxRrKzy3n/Xw6iclOhFbEtQvgTKn13eVU33DaxH6DLG9xZ9CNDMqiuUNjEAbxykJ
2AUrnI4+4pfh/EkeEFdyf+zfT5y+OTvuTCU238E3H11z7GkldbX6qviubQYX74qUHQHkdfSISsMK
ZfRLE7C3kbKaVkL3kOeQaeYICPu1EfF3qjgPx/zJKL+YulA6YVK0AqFTDzhzwac64f4cEVl6H6Ry
JHE2ubO2Eb6wqkWwu4UVITsoMVMVOyreus4LJnral4urR7liMG+qw9dt+5kTfqW0a5vnGGW5B9H1
jvX3ox1HrsQizF15MOiF1sqzegjAlT89hQD764Xd5SQjg4debM+Ce5dfPOsk9ZLsOem+/tRcHW0J
9kYfLcAeWAGr0BcWAU7TNSrf+m5qMpOrY/QgZNh8q0WGT59URmXMyDqQI2ZDGrD+GjoyoYNISgop
5z6xTxguOolgbMXv+tfzY4IJj0Wq1Nw+x65O3z4PPgox90lW5u/IGyPzyDrcHVzn0KLYexe0un61
Vv/kmHVqvG8rdu7rk9o06uy9EKBSTBhkJgf87HSF2yF6wOSOtslpxu0yWl/ZOWzm0/+hrbWCIRVj
/QG0rg1AtVMJRalMB3p2WSwcH/aL60mQurws8I1ac+hvW1gdwwWJNSCmiu298gRSnFJQulgJMlhX
AbBq09qNGqtyIgKAFfkUU5cS0tNhxGsS8xmORVLkXwszpXbOhehiZUGl//xdJz6PHJaR+5xkPa1S
yZoxSOVMo3nOQdXskIHxfJldPbY3wPrD7OhvTxNMhbkBKzpdKfK9jQgF1vji7QxZk0wRpFo9rPu2
QCO5cdfz2zkJbU3GBgFie2v4AubpjOl9jKXV3eopEyROCE4gwtuycF1ia0qq12x7wjbOfc82u0zj
JIJN2igvoLhPsEZWO10AaHoqW6IvtCv459DEwgCpsiKZB0rN6oeynK6v+vOgVHzWm5JAo9j8jayR
RMIJIrSZQr5cH5h7FJdvaPTgL0pWxp7iJIOKf5WjyJaP0xlnrvrgfA2Dl3/hcYpu234l4cORSG2J
6El6wh9VcTcd+F2BN2ggKvtZrV0P/Bp+XVr/X7nbyPo42RbrIplPk0gYzoDl1wIoT9XjOLwLUaGn
lNqbcu9iURl+Fq4ksJCYrX+JXQJ94XNzyrtMCufYooy0dW8MV9idJuK6EHqtyFB9BDDBwzYXSEHa
3R7eXeFok4n8gznuwC+iFmgAyXPWCvg9/xQ/TJM+1fiDE82JFhM7LMu1FcxvyJPYksunhHNTT4mo
4b82Zepl+tfYtPNo9lhmm34SPf+uFc7P8eO+llYBe6cs7I4TQ+jGPYiGtOOhjk3SqZegYYZPEMsV
HEuHE/S4oV6a2bbGbrpk4MD7HrQjXMuiS9sew2BVLuFfGAKbcTYAmbadOtgm/MHe5GRHUKu5Gy+Z
ClHTpRMB5uO8Ljz1ZtvImrxTqg4siEyXMxeZuh8ITo3RtBpdpQylMn0c12g3GzKswuxLxQew5F/2
8G0xOjKmRD380e6S4+/YPSHQEBnKQVDznZmPDCNX2YVz21+U3o5pmjG1s+wUX1N4gAOheypip32A
JZoNqlkfbVdRGReU3wmGlOfZR+KS6AcRw3X8UfDN6N8N+YY9XpPerucTX6GJNJQtTIO808/VpVdc
jaeACZxeau+U9yMgWZfzSwZ6WmKpDPnmKtyO59cYVtSchyu+7UmrkF5NZN7zZJluSNYJI3H5W7jJ
V9GrPmbZY6j5PBKwegZZZIjnapeCCT9nEI1M/lN71iYXXwpkfOMWeMd785TLtcSS0drMtPQVvF2g
vrv1PVEOodGiLShBlrInVmv8hQA1H+U0pPnuJh23Y5P20Hddcdo3GUq7gIMoWnJiDcPeMZBb4q0H
ifavEbaeieO1kSbqkFium61W2CQp3z1/6YR96+Bp7598RHVMQrLCJ0+gihSrkBZ26iq2MS+BoHQR
DRLEEZvFVfjhz+ylUQikiohGvE0YiIbZmFp0DTUpAqYDB22NnDN8YOtPKyZ5dBQKSZvxR/gTb7B5
7g+bqPgz1+mYZk+aPm5uGSZA5S35zOfAhbg1wRpQYb5n5kfPqeeOGW4QaWRcKl9lsWQ0g8AuWGp9
AaROv4kpSdB4IorI8MCZXz7DEzuXTsprpfJ2F/bwfe47xeBglY1zLsIMCc+/6F070kCy6yd1KZw4
LzperzGpXevSzvuwJP2Yz+0STeJFwHBJlrsy/hVN57qZFVFJvQ0GiEeP1L22suKKUcsNVNy5o9a5
VboJLoxv+K7MDThgVW7rVdo8lsAHJtfXCJeytbooPiK6z3f4Km9dq3knF98AFXyEjWxtA0SfLzQ5
TxVS8NoJkPvK7Yqe7l3l6UHhPCrNzrXp9env5qgQsL435cvQ8z37cAURv8x43uwilvSdL99Hmhix
SBwP/DSJTKiiwxdeSmrU3yXihLlmz1ePRTF0xEwtm5VRmCAIl+UXNt2fykUzOEnXWfeG4TmB8zZ7
LlIxMgq68bD1mxSXM8UoIC6HEpdWCFVQ2LQ1zrl7c9U7CJe0RgtyQEkxPuBc6BjlxJRDlvrS70Cc
BUv78/JcpNOarspAX7P41ilxAfxpXz5GiYka0E7k63v3PGFlCKWeaylfPS+OwVNC7vEx0Fd1Is7i
J3s+nP9QNaBrIwElThj3HJ1eJLZIasB4jqdfCkVJdmeb/qUd1/o8I5ihy9EgvQvSMVsxq2qR0Wtm
y/oVuoT+gvXlOwa/UwZE8Gc/e5no92Sg1Q2y7Nv4mOD9qImWVXZHWTTkKejZuOhgooE4k3bXTxrl
NxySx3OVaagbPAjo2hQAin7ihchb6kh8TbcXJzwAqJlLjdvUJBCwebRmJqwseJ8S+5524kUuGNwY
ynbpDuilID9NMBkbreBsdoIYy9S1KDWv1TqkWtC1BEJ5Ho/B9DzOub0SO03INoYjaylL9Ekd93Jv
tjmDLmnSHHWyPIuzWSlmVE2pZOgh3glecGyyPfj8/0dbx/IfLb5mwkzqgx31AH9fdjtf0dEWnP4N
HFdOJagUAJaPD0FOU3FqadrJqLH2+9spUBMkbNBsVR1FNYzwhUxu/RmWH7BVihTAlQH6Zi2qysAD
VD0PJ9lHTSC7i1zgEXbpRbCxj3p5J9ItTzrs4WTivb/itJp7X7lHZrVhH88RnbVuOhsegLih4CnA
F+v8NiWYs18o4TDcFFnMTzgOO28oiLuflbXRonOEBjUSh2wyi0+KeWDFB4Sle3m4xVeGq/pCcFgQ
RPxIN42ivJRmQ0LPnn6+6tjukXUaRwJu71xwE40XdbsCLdy5e6Gx1fbHJbvLBne6oV5lQu2bBwA+
+sftmhGeuEVApzrDgKhKx4kCf5d36JtAvWE7kX6NLjslZRGWNpYg2pGQTCJeUQe5GD0Rm/W5gKwp
vtiDBsai+4H+UcTdUqRFT+70w4fyStTrygmVUf3+nJ9p5pSkrHs9CF/6da4T6ojDIdTK6YO4ipzD
xtZRKNNPzjgVgW0wjHx4U3oSigrdlaJalo90dWh+nlZRNtykYmraUEw6yuZYJtdMi68AL+6/tPO9
C33LTLxc4MJNSn2WjDOF+KGBDgD2oNdrfFsAUyJjuJMQCBSV2YkKGAqhBRFwe+HOZeHm2p4B8WsT
QJAoDEzD7aWgf6a1aoT0h2M/Qm2TppvaAfFJnuJ+P24YxfPvCj3XbQ7NklBTSSICuo+z3b3J/Ecf
fgUY+qv0+FYPbKdHC9EDVLCljKmnWXduOR+HqRNt5lyaADN43eseZwXQemG19bN46eiv3qilIiem
9rWMnuZKZQpL1imWDWUuSLYD67KuliF7UpCHaXFg3ra49p/ixy7Zz1TbwqMCwv/x12jdZeFYBnhi
ESEm+Z1x7DQib9kvx9M8Yr7MpFQiD3caE3NCuCCUdue7B6xRSYXuQSiAmd5kcsE6oExGo7L289zf
6LTDhs2lo/KlhIWAJxpGFA2tqz1DLYbmrrVLSmMXyuEhc77o8c7JUJTGe0uVey3Ur/kdntXFVKzq
5sIRrjgU85ZWeH6KjMzQMxwl+04Vq6NxH5CWhUG2D/H+NZuVydi8atZPaQPebEYwWphFhhfKxP/E
EcPyKKqUayQP8hoHI/oNgmagx/B27Xd0c1GcDSTpCnf1xlVvxeQ84PgzLxCmCFlTxRF1zpOFZMOQ
+AhBPLJRKiBiN9mO1oyIQdOvo/sy6Epz6ABna+ezgVKRGbeqpB/xgouzh1r5JgJiWbO7mYPwlqH9
IgVFcA6lAJXJsGdI09jfdSkC0RnE2OyseiAKeOjw+aXRhNjHl5MvhXYLc8vQIPYhtU2Vja0LizBv
40T2zWjLkN1Tbvzt25uuRWmK5ain0FEILTJYidTsJ+E2CubFarsM7xDcOPsx670pOx0CsX32Vz4i
gyINB34jB/pIxGM5o+/9wDG9wIg1Jz205Xz9wtM0hV9MgB21a7uWhOn/mAXixeRCGadHR7eXzZsv
gajCQUNq6ONp4N0X7rzy3/FVsxGxwb2oYl/AuO4wkn+KTnq5NshP5y4pp7o+2q8GWNNMgjAaTUVh
DUf47CYPcpyDnKlur1GNOnGwhmj/3BYZn/Vun/lNi0weEBFdjmPcre4JY1iaTS7NayCdAFCkhh5K
e4AKcPUmCno6bAraUcUGL8KppAYzB0r4/8EMyjJq/LYQQ/+p+oNYVPh5JZLxvFJ3Jf0h1LyeT1BZ
2KVbHhin5VZdMFvcxycdzAb4Y8xywxgMh6uICf9YaftNXCdxuFavk6D4seJ0pMNw2tgoKoUiEW7k
RADwJ0jAim+9QpO3t7zH79YZwHsILbVdZiYUDLOVmQIfD73AAT4zFdGpxM4S5ycLf7qcA4uWiRrz
2DiMVTutvaDSf8gm+EOiA+8ddTfp5Qyl935b3RMiGJHkBP0Xmy+mww7796LUnG63qcol91bpUWVY
77Mh4rVQrsNZRUigFgJhb7Vx9ImJ7eWP09WkpEglaj+TQQPESIeOJpowCQhqX5iQPtSFyr5p/9fF
scaUOWwit30gajgjkfnKdLKo2CqlwVtRUr5wuATZiOjXU2WbL+b/OiDAS5z6K290Hz8DDOFo1e+z
djegyLa/9ku/OgIiEotD9V5GzVtURjeC3MgXuPvcEAuxkj+IZn+o5uyuZE7eoyHHeo8TmqTeReh0
uloBAQMRh1HJbcRQoiEL9/J/zF5ags5P2DGwzfO/VqWeXvxXmWZqIgzmVTvXD+5WPGCeMkpJc/X4
bv9xQxBssISsSOqECnMVFgLloDI1PBWzErPBu7+MS1hTE3GLJ0uVONr4P+f6HBWplq9YW5hwuO3t
kAjv0Gr86lkcwSsIr5xIr+ElpDYIerd0C5jF8XPYlc7tX3peLhfOr7Z1KRDo0Q8p0eTKkid03yqJ
Aw3Soz/RcmWxq6NZKL+rh9ktbf9yCjM+N4XzwlNFxH1PVej/z2zY4xoYxWgrIQINf3LS7cl3VkUa
fIF05vbZx+EUVMycgGST0OUOR/Sxo55xLDx8oIZ90cqZzfGEdBGFU3hYUizuFYXj0BbI7iTKrzLK
jLQp/CxCa+XJR6B94gE/2+s61leCgAztIO0ed5zQ5ek68K8TlzSMd0QZx9CtjVYmFEpbb/svHhIc
ITvxQDNbYiJoXUy3CUXNa7SrxyxKZDidNqPe8L9VZIi7H7d4lpB768FxmyNCevk8dRxDdITJhPZ8
Y5ocAux3Hdo8nSea7wEJJPWAgMSknEQviyD4dYUuj08hsy+lnbEcslrCyp4HlKCBgWYvJrX7w7Nc
mFzJ/1ixCk8X3CGXQY55QiOu28yn/SrPcYgAMSmALCgHasr7MNw5BdDbV3cTBvjcF0IhRIDQqa/C
orVqdorKBcMeVcAxBu9FIMEdJT4xxODboS3bCRca4jRpGPjeNRS3/RZ2V5YazsEMp0kgaa7U7kB3
OLIo6lIqWJE3wWz6V9D8KFxaVAwkzlLSrKmlU6VqWiw595+vXlF2zPU78fx82VftoS5kLoNHV97I
edf/Bpkf9R1NIkyjn/QVkq6RzeUHj3Lwa2H5q35OEyMBfohm7DkiZSJ0cfO+TgmEx8R4diYcwLCQ
0Vhkbt4OdKRr+eUOtD59D/D7Vc8pUcZc7WFnJzT7Z23ODTUn7X48MnWnF6qHSitwVpYBKm3Y9bnB
gSwVXN9C8PtSUrP9XsZGSZbzWOPfHqGCBWiZAwWVIxvPO5VLsDdENR4kguO1jTa+2gTu/4ZMkOOT
B3eFnEKmta4Bsah3cMUut42e3f0EAAgmB5ByFTWI/SDgRjLxa0xKuxQxeexWpV0OPkPeov8/MLC5
3lOBYGHwaKACsVwNcTS1d8kA7pNSBvbGuoNwYkNCB9nxcw7uP3+rP7K/ETen5tgBMAxs+dvyej09
mO1ArsxNCGHNPk+0LpslEcu8eGd5mLLo6+JYx7CYweVbmteDPIPmxrfzNypyTsrWFjE+wtH3FHcR
srWJ7pBdDa17Pg2Y/izjOZL6tJ/PeO+nMdmlzZJVGQ/d5gKruEOZUW/v/KqjnCsvqawUrer0DGO9
aTgEAHz8rPEktBp23v7OrVLAeuuxn1HKXm0p+vWCt39KNYYFw2z1j3VTG9TEEW6spxIo5JUKL+ay
PbNNYA7beC/b9QcjInje6crkU0GoSnu+zg9Yswxe07TGrwa79wk8kJ61Q75ss5w79YIJX3OvD1hv
g9MQGokJ+EUUS+fcLNMiH+310TBe9LiKK89wd5M1t7BuBy+7wbluNAoVXw8ke44mClm9fJc6o59Q
eEMNWS2uFGfUeXMNQh6WYz6JGLeHl99I7uedcJTYW3cyJE83NU5YTV3n30vyKnmaMpjQClyaJxD/
l7jzzQ9Xkq8H/3rjYKmxJWmlFl2mdbivGVNRHPWt6GEZ3QOz4BkshhLe11vcrYHsulLR7znLnZ96
YyIM5313sdYgpsYeSbpuR1KLKb11J+Ry7gsGq/s/KZD1gzJHPQhk600fiO5rTDPcxsO5z4edIsU2
3nLYED5A4MXQK+h2Dng2tdGh5zJS6r5p4Yr5M4Oeh8SweO2PHK2tyPIrBJcdT4uud/4deRUtX+ji
ZKbVeIKYwfHB+5hMHXEdQb7a3TcBrNr0kb+oqSsA7kJ6GOup2WoUt6YcKUOxz5jJU2mrVa5L17ui
98v6DXgiKrfQ2eainScNcXlkKoSNnXCUhV5buBkX6EAKHdgT4HyAbKSOUbxFW1DCLU/8irX5PaJa
EhY0+JQi+yOT4aahTNxeAUGKlHnmQJ08zE9iOQMfOxxhbg2c+es/2FJyDEnIAuHEBvtcB016Wlrj
zJGe7gI9b0vZLXNlDxYkkjjNn0yH2T3WnfijaMwXt62LaIrtZ/kQSZY/eEm2FDmZr4OPcvW3wDCe
VvptL+nhOqb22yc3wv8Geq70/ZIfq97iKx3G42BsdMMDp+LOgou7wx17Aqb/mr3iAqhPHUi6P/uv
TMoZMMwBaSsV9Mpsa4gpp99oHq0We6WSip4u5k5+/SLEcNP4tyvRnnwlXpcR7SI1tt2BMVDt0FPV
9nvYHF1VWUryD+acxV13G2hnAe/7zaWy88lyJ48V7xjhC9jzZuQT/bld0WgMTtnQVNoTBuynvMwD
vFZ/W6ArKpvTldbYBrBMEKjpiL0/m1x/L0ZFrg35wRy1IEitj8dVTmAJUgXC9w2hji081egvq1Z1
kbMR7FnMX90jmyIcPs3nzJBCrReinO7fIlUJoDOEewDB/A1G1oOJ4W0GH6iSqW1McRssKelmCZq3
kHteOQBvo/KJ2ZNV8B2voMPxDk0e7T4F11HZM3wIjYuwRsfMhh2nW54f6VeITUKrBi8wmPinbEda
tJPSvu8/nPrk8N7SnXu66kqvVFo7H2V+VZ5jDR4WPIFvUFqgLNRTr0eLmpWf+0aYF/s/6osOXZT/
0kAewx4q8bS299qKRN62W/49yuip2B7gkoTZaW0nLNjYYSU+9TMHamSiIT74ZFsGmOXwUh0bCS1y
RF1f/k553coWL+NFFWLLDzjSqXvjrhBjX4LIPjEPdbzP0iLuVC0rkU18QCaKS/D3Q59vhqH2LaD5
N/wi+zfx/1Gh7TW5HfIReY1qfn2x+elnqZ6rxdZHPb/2agN33UwA8/u7+q/lhXCTrp8Ql+vKE3gs
twscP3Ryxhn1DhQd3IHpvsg2ditCuDsP3xm7UJcYArmBYLKKSdA4e6FVc1utmlO1uu/DWIP0oNJ1
hilYqMEKLXSCJLr8oyi5Ai8g1XlAqEWZfb4aBccF76z5B5O2VVgjULaUBa6zPCdGAdcEzVg38TF2
9NMgayjCNm8tIyfkKtB+QvMq8wrfCxKpnDGGrfxsoyLyQ8D7NgKwlTksy3uYU5BQ5WtHhufckwsd
XU1E6iwFtiGMWeYr6/XK8BPHFJcyvjCZRLKikACqFXdhXr/mSgxtbc7PkPL62L5bc+FbzJF4Hs+G
W1ikzxAw/2tMCicw+nvsjIEYwztXHQCSK86I/W9xldOBj/ie+qZnBpWP9kgtoO957nFtzPxuBEOR
KyGF4fI0oBMvGxC9slkX2XKFGxhzmWg5DefMBduS8vcXAB0D4H+iDhLU/LvdQdrnRrTEjyrx2CDk
XiJyeMNCNMUo4BPnhm9438hr8mmS/pb55H6oJGDq1Em12UWxUnfWOn8+r+E9ofA/cPBWcVlpCjKN
Q40A3zGmGfWgmDqPR20EyuwzBbctahUcuB+CD9JoHeOAivPWjRFNXVyZbPslQaAAuFUHvBc0zp7K
xWwk8gXGSIrDmJsfhGurFBrpTMFxY9W7P5J2lqbKa3vb9y2g3Hl86mvsXKh6ykY5SD2FkzrDUyCX
1Q+WBbPKLIGVtWmxJZC3SBh3nFniiaLlf+pkznnIxxcaI+lanp2OgRZZ0ZYEyradVRNhePUsOWNZ
xncp72ePQrgYSEgQifqVUMhP8tCXoKF5rMkOIFOY+Z3L+EG/FPm1/UvU9GLrh7w2VDY8CAtJWvTe
D/7x63MgFu4fMkch1e6zfwkVK7DF4lLIXOJcVheoqkwfGsTonzXe33eP3/v/MCrLZYdmCkNgK0NC
UNvBe5V/t9ll1jvPvzd7yKkYo7gsKO3VM1KfGDjTKISyofZAn4sQ3ToJs39G6My+yhhdqrChbBXw
KeDXQ18QpagRCkq0SFYDKh64wxH2YmI1gJZIE2y/vaGU1qmYBmhFRVJ1lSYIBIdrHxAPiAbX23pQ
ExbSaXeawBGVg8Ra/DsaQZfMYbpKQ8tcoaK90PCCiCjKkRtBit1EWmaQmOyu3H1C69TOjnZuzf8H
dGisQXqd3IFQ3E0fQZWvPmbzBuPPv84gNRB125C0k6H/CIOVfZEXj9WdDWPu4a2NlnxnklznZVo+
Td+M78KrpuwjOAkmAyuVCUuzOa0nZ7R+5XMF5f+GRkDjMKjRC/JGisACeEbVjSZ5CmuYclOP9Xn8
AEBGsLKILSgNL5LCA6IOtFKJK5FMWm9APOGun6BkhGUJ2OGwPtCPBt+Cp8gJ9nIVq9XRTaeEJAYZ
xIYNOzpH8PLewFpgsh4tzq7PplsAkjmMPOmgHZlgMn5RW8tJWAgojQQZ2GkYHPi4six5Q71FWI9s
Hl/3iQ3F+hJ5aOLF4Ey/ahhoR0FTgceQWv2y6q6VN7fboU1SL2Nb9aoJpRqO4iE7soras3uCLizs
WncdqythyMbRtuXgZ80Rphup70BNcf4YerDomLNn6DoiLRnlD4xFjmEiSGuklqn78B5sojUwq9p4
PhbWvO6TekmwU5wmOYW4rJitCdoDzV82jZan1gLk8wcu1owMGlbI5V3EAp9quSQq83UD6M6Jh5Vf
xY9Zm3a5hNKxGGiAtXv3RRg/zJ5XeXJCt4RQ1qx5e8TiAIix+b2BwCdaI7Jnq+CN02FnkjJV+9OM
8H1EngTBe42XIfeBJNKqJTXcjVVsn6MwNL8csRidcJ+mSCAtN1hWCsX9EcOO2c3nLrzI7WFF+sAc
JCVyZZ7NhmApZpq+lr2+sN5xKi+2A9aQlhZH45X/WL9qUlUwAxS/0NHdigug3K8qDOiOezIG70Tb
G+qa6mHzW9ZapGiBFNNsLVCU4AeRP3y4vVrcZ6ZL85RZnawCfPLFeeVfvyjjwmcBZE/4TwfKgrxx
kQUU47u6pm6xx8dpnhTF1zOvctieLbmGgkKQIs/tJ01vh3s778/x2cGnn84OC1eMtl21L873Ef1s
VzWG8yBxvvMGUKLs9o/yDy4zDsvUs3zVIn3sHCInq0Gpu9U8rJo46NAnTvt6GBvmS89/blNOlX/Q
GBcbBoq+nQsrV5FbuarR4bPhfEZ9BmnvO7gNzLTv/mlpRxeWM5RmzU4qVIM4PEbO0eqAnzvc9J43
Yq/6OkuBTkkhDY8XxvPD5JbaL2DfB5YvOA0Ao2U6UTa8HHaUGGomd47djMRr/dsiuk4H4/dCmnQp
A56WvkOwjNqTqk5uso5INMAbnIoeGUzF6VytBpyqdvl8HTyKQBbfyG/kmgGJOXgCiDhrMxKab7/B
z0fu8pE7ulVVfu13PxhwQviLeejHV9Ze2a1iWQa5nwL20lhWPxKLOQASyH+QLNytY2AHGjbHMDvn
csFryk6v1AmEx+38OaIbLjrVWVZbNsowxzjO67EmU/+EWfSYi+L05Na+9P0HE9UKbyUn6Y2YeAfI
soW8j8o9cigF096pX2+H2cuWmTBLKNYHyZUAUrTL5CTlKseoYfa4Q4fTIcpjVdRciXNG+Vv5PfQB
/MS8LvydtD0y7C5HVO1FO9UEv/rp+1VJeJf5ilK1hyYR3ZrhWx4wy4EPZiVbiKCsLoWUCmBZadOh
fW5Bc4GJmnyFGeKRE7C5lPcmWyUx9MUjHA5Edxr9Cg1cVs9QZ6nbgwWJ3f3+BzQSl07PKNsc86ut
V9VF56+4BsfigdGt4+7B7Y5roElzZAePxrDPsJxmsg8wXuHIKiSy+aZWe1rG3ZhMicWiZQDpmyK9
CCCaMOkoueMGqcoxVHoE6A7B+3pWdf5stkh+oRNv31WK3Pm+26y/fipGbbJ3Dv9urD2i2gwwH3qy
ggUPVLkCTr7PPN3tYEABTSyOAt0HHsT/uLWtyzw6ivnt6ICtQcig8Q75tC7l0zmAMlOlqO242CNs
YZlw5Uqk4hmUIi6K3WZsIrUATI1t4+jANHqGi18T5AVhUtZ5R2RwCyVB9cGKBUa5phOiLt54rI2i
bx4VAQGv5vugtUtDfN4D6WClpre7eRFkIBSmGiqV8bk6OApmPT2B4dO7NT8ovan4xrcPpvZFvWxV
ioVuR+wZ5vF7Hd68Z0Y4UhcfCeCyhmoqBuBd/CTiM4m2jo3p1IsE10IL27X5XSRf3lP0ancTcYtB
3ezOD3BRbYAk2lSDbWk3M2VNYpTl9Gs8XdOoOXOOevILLYQsd3LS54qLEsf0fYhLd9SgT3MgoX0J
gL3BOT+iTnNY4/H3eqZ4xabAqqcX20WUu5P+C2a+UwKqHfz7Kk6suVxDaJ06G/uqOSha0Y4WrdeJ
8BOv8IGdrqcwjMDnR34f/275zHM4GFBe8SRHsqqSHBFQNhlM2tLDyglmhLhakCbspfs8ObQUU8IO
u+KIbvMhzzYYRSjpyZyhmiPrVTwG3oGswLOuMAm0NzUQaQzRcwZjc6Oj0H5wRvLki9lxhlL4WOk4
Aq34HZK+P+L7tT48y3VtxBewK1X0cl9ZZVHlQ/II+A11IO7OiIrPPyKO2aU41dRjeH/s68h4vbFr
2umSDVnugtWKE2quf2rdfP6ilZCjw63e8XeprlT4GUr6mH1F+LRlPMDJygq04RRvTPY3jHzIx7NO
LrYdp+s6193GpVd+CR85Cm5u8x9uBoJVrBc6zKY0aO6khkJljVLkKnoccMPnaKSDT0wD5fCUiz6C
BL0IFJYc/GToB63WTKxzR/ue0t712VnjaZxMFqfO0CcRfXRSZD+tJopuVuS3w7HAd9Iduh5sxDvo
RBm6+3mN10fBEl5l/7bGjxp67LAhHm3KsFlre/9edP/lUaWWySwvQg//JLI8bhLsBuoMulAFRCEl
qrNAv8NVnSoRgA+JDQYJIW7zB+RkGhlX78N7yD9q/VzisR/fBqfrHnCnVB3pj9Yx21FY2C0KInkS
G4ihrsg+dutJ1y5S3de+DRKRwlIbe8lOmaOnKvzBLFTPvWXhPKcPCD7WB1fkRzPOVVxCvZeZtWat
GTVMLhGw+Ru2D138lC+ik5qvCrk273TivrXXWGhkbxVcwmD/Qori165Iv828Dix2eLVSLMGOBcqN
cTOsoCrZwucsKAsScuOBvop71j0ZQWxW5hF3lh9OofnfkJN79GjDfKlX+B7gv4THn9JxjXYwzWiF
ZVuxVHz9xeTLs/W9Gqk5EhtWU7UXsuuDEtETX0S8Ydnl6c+Xhg1uZAAGZDTErLkKsBHkuFJR8//P
tl9cj+4rjzQsGK1BFi5KneoW2NzA2O+A++/7Zt2aUDuqMEg8EFOpFxPo2dSFKGjS9XP4bk/cdVRu
IwJ3yb90vW5AbHq1gkcPBoXqwjns5TyVyPOywwrQl4lccaooeYR2WA13o9Kdc7e5FdN2IVnSmxhe
Afe+paeJeuXYjNnLrS6C9NbfclfBZ9i/Rhv8m72Ps+sBvL0nAGG+Pl5XC5RzxHQE80/AtXSkIBzy
+C3neBgFnEDjt3UI9d8eep9r+dOcVKfIa/JM8383UcermmqlGH1AtuIG3BuZsl6wUHJwy0hqZoYk
9RW00wRorAy2+Cuqp7DzQo0w38ZOlr+Erq/pdgUw137gjTa48YcPgPsP6F2a5aHJCEP+PgkMzG/8
Ne68jkwBFBDppOQsNOSK4FOkZTce44vIqemCQwQRednT5T2wcemsQVGDWW5GS+9vf0dwT1my3btO
2OzlEmjVDbCmhIXw8DwS1K7hugafE5/BpqyNpEtMGKXIGghzia2CfGu0FtR7oyZ8+tfrmEI9VnKP
SpkU4spBUx2ruF9bkKRU6ZF74opShJLcYGVeBeeI40bwCMerxkgr8V2qjs7VGBL8CABF/i8mNkzM
tHKPp0vVk6TlwRtLTK+M9ClYCR6HsglY0CMlm0j5xDE62hnemZknrAvb5e91L0KergT/yhfduixc
8ToHQwMNabdua2tnVLiviZj/toRlHvc1h0BoOwo+s/TRpY4mTubm1nB1AWdVEQ0FdkqfIEoJQeOH
aiEeQ3k72Lo5okbUCuHQKLq66w49CNIdFGugxsqeK7vFGAQKGnJtZL909WA4ge+X7K/MSR8/AyN/
2QVLpJQTbxkMSRGhDXs1iMOQ72/eoQRPa3akvpwKQ5hlW2oDIltPLKGOgefA2tTxoo/t1LNqyXim
dYQtyykMVn7T1qbWT0PBhEY4tcfXGpDDYBjHyabKLgFUOcYTu/g1p2ODrM5MXXuQsc54vVG84oXC
s9XufxueHlP6hDuhLX16ggYgdx6fJz6c3+mew4xS1ZTyuVNjWacTyL1GsJQkIWWnUJ+b0mqGjHeL
qggyiKNx6TQR1x0oak9l1JXpjFC2/B73/F6d7RxQMaxNxLsH51gFI/VI4a2CuJnq203gwGGjFGdG
kS+VUWb7gFkw1TB4Eqwmp72kSQqbg9+p1zr1nwEX/5IcVpxYUsn0EVUtjaN4tHiVMJz8+UHlwD2Y
SuGx7oaUItb7Id6vi0BXuedqwqh2LwTqS8gDbjShPwNWoupmt003hUYRjhGSbOYw+6AA2zakIIY6
p4WT/lp7haz5jd7YhFbpHVxGUoEqiX8tge0U9gZMVs82u2TgvfVq7gOnAfvvMHS6k38mN0O2TBGO
QzwIgLI9aw+2ekBXrHEDuWN3qOIlIrkdFucvUabnQb03kXUKJaXDL2hMFZDacBKxLea5sU0c5+Um
SubouGxgBYquT8wdIHVTPc0l7bHiPY1vV7A/xfwBZI0camNAgzUacgcr9nZGMefIG3JeCuWr306J
oWwcLK9hjF/1DRDCzBj9GOFD5pI98VCNZBfsjDeCYXTUuiQLpxSNdeYpr0e2eSCoTsuP0t99TjWz
TcbzjFMCbJhVYIbxqel79invQlIP+abYhl1y0wN0TbQ7yseZ8ABr7BFneFBIb3YAo4XQdn0YEmFn
9bGa/cdXo3S6V25mZvmfG/7jxxOLScuWEL3Jv5ATb+3HURgcg8LOPANZX+m816Fa68Hb2Zfvb9dc
e0J0SSFm4Y5QkFD+YqTnYmmO9iC0pOxUDD3L2adllwavCKENlK9xJhVeMpEE9qSBjOKt0OBLv+lQ
SWmX3NoBx4xiE2eOMvzbgF201k+2TtKXFDFYvHUtOMrmSwvwVz44/wGHTdVBDvxb4CwSlgQqkKyr
Lh66QCTLW+oLvcrT6+bxfZpv+rhzbm4UWxwO+OKtvmwSBzvxSn2pHM3pC9B1Jg0GAoqJcf2MlBLD
2FzcSGh3ZIg7Yg4A50nZ+9Z8Zu5DnRcHxEMGsqBKr2jP+gWs1QVpV+/AuzHhbbSe6+xAFiveSBCd
+jVLTw3ZTg1085P8Q1xmPbig4toZyjmbjxSemfzsQE9Ztne+NzHIK9QTa7XNlV6VL9TS031wqons
clRoqMP0paGURa0nFY+rp5kEU6hcV5BMt9mWtyVFlvnQ/8ApIjzvUXfeuqbcvM4ap2cSFWLJIofY
kH6IMym39bBNtO4x4TYX3yi0+3O3UD4qNtmrHUsnVfgJfNvUG9GdW//kYm7cfzRAmOtasihZQgHH
zsIVQcMYveEelkHdVN8gwRtwFK3q4t/3LshpPhW1Q89bKlAVJYvN5gZeMx8uQd7t7gsELhByatP1
lra9ZagxmMQtD4PvvuAf+HGa1+LFPefSpy2MUm0MHwH75zALrBIZD6hwsFz4A478ijotSPCGnsAh
wdeCXDJcWmRJG1ihBxuHJfoP9JQWgXjZ+qEw3HxWJ7J5G5lKAE/NX9xjXoVyJcsoMRpfQw57saoJ
BrJW0KTaE11/JqjUssQmIZkQHTyVBro+Gx8+Ag+LKo95fvaDdhnoY8UoieMjrlQrss1M1d5JJ0BE
BtGlq4yvb4evDM2Up0r3lHS39Enr5Yj07vSMJvPcG4/5ggoCnx0RV59jj7oiQdAesIi31itNPW4h
bCAyZXN1Ov29D8fe6bM743OFcjwWZuxQhML5tMj6YN6pUdhYnoct/s6SAxuPpyRF4tGRnFi2kKFT
7Y/9uCXVKtpvtU6D8hRZbhB9CUs6rezNGWCoxgi6t2nW3dVGbHAYkZAy7g/ymil9QCskJBoM1uPB
aLdkd9Naz14t0VkEUK/HdDwIGdcphu8Gi531K8n3B7AkREnjUkR/sBxWD1yh04ZLXz5v8vi2ZmQL
6baY/ZpV0JVBdVN8atf/iHq5f1UyBPyBfVEnLyHABYscnDZeJWaN8W/X41sUymNd7U6EzUC+i4Nc
WF3nw87XEZVed7mHA7f0IOhZIAqmqB8MKnGvus+Ma/sC2Pt2DUikDotfaAgz7saF7RJHmURLbKCU
Hm3UbtkXebjp84/QmJ6Alecq6XXMC3qDxrNBS9OajshU5rE7zlORlhuD9iBXJz8ABHZwCjT0nD+Y
kyHrtNy/Y6zEz/S3w0OiswBR7fQsAVF1F8RKzRUrezConUZVSO6Vztb4PktalBJXD5BknMojiJyI
PJR626kRu+EwUFRypo37tV4fNySOv/0H7NX9UO4thCs7vmRwoGCbqmlvqqh6k6jxvogBrOQ2Mo34
d5lk3c2Xjs+T3J1DYBdv3gCwthhBLemWYVI9P6u5vUZnoFn+NiZ1x8MPWwEA5CfrfgAfMTHhIdMQ
TmP/7tbb34C0dyr0jGY2HyvDh8/7y0xKBJOxKGqIYGVQxh1KQbpFqifgLO8j0wNYH+AUsXQmg3QA
e5lC2Gr3mDxA8Y1rDzW1ek9iBqTHWC5jrKUvyrZbHKwmeGCENFHnr5Xq/jUjJyPwuw7d9sKndPJD
ZR8da4t9oC6CNyEUcxaB5zG+N8jbHN8S5DmUkzaKNOxEW3VXbI3CcvxFJW4Hklfwe7DCcvKKuFRf
0Cga9BpJn4mtapSCv3h7kZ9TCGN33bBDS/CPLWFZ9Z5ut8eb24XvExU5ZB1m4de/4IdlYLH2UcbB
5X1rLpyjmiCExnOMhqyLEidMQkY5UkOOhEiZus61l0NXl0PIiz0pCQ7dUjaaeefuPNNDcqcWvsEI
nWxpx9n72Vnjhrfn9au/MRrRy6eOsx/vbZpEvDI7pGXfBNkUyZg5dv2L877iCcKnNFfMa6OqGIQP
HgQOB74ysR2l28dxKxvXntznLjnh0eufhR1in0ItESNFNZXBWNGAgyq4RZWVcQG3UbvSVyjc/9Pc
2qLdlfHnlIlKDCD4clvm+hKrz9w4r8N7ytud7u58yTscFAtqqMWksd8He++bX+KjRNMD+UpTeCVB
OMH+kXFKi7po7j9qfX94rIvIKSkuX1CNoiBUktBOsxKGLjMJddwSpqPS046NixwzBZkpfhOyNvfQ
DdvW39rEKpBtS6bwZiPRdLLzfpE5AZwiJxMnn3IeTp8t1e1SOFh4NE+QeTp0IbK4tOarAWKjVN8L
w7y9HzgJQzj0BGyr1yLG7XkLFA4tyX3hDfWuaXYIy3WkQL0PtijqxY2waKtRvzsWyFw2t1s5SpM2
z9MC97GBy+c+uLB1A1I1VSr1zCdPEBkE6zAk0c+VinxoaIs0sDxK4oGE/olMb3YcF+n02p1vgOYA
fkyuRk/6amRW2BSqy0+4XQLSxIKADSiacTVeQvMR07kqVkDJvfE5n3v0ufRZu2DjnDpm5wMeRII0
yMmhbhP/ioUYaX3AgNtQSXi/FZuJrJdDp75nGzoarB8q38vnVbdDcfYlsw/4HyQzmE7fLH4f2AHN
JTfwQsBe8uMM5wVH+KnT0STh4KmkD3cgtHBEvQ6Anjz9Nh2NP/WuCdwbowAZBwosjxW3bKGkBavl
QmdKolm9P1Y8doZVji74FeULVyJTS3pCuQ5IHTAwsdTuQXILeHvJNH20mwlyejcdWJgklrNpDQG3
CmSLVPboE7afT/ojuHZRQgsIcTKCBkoCsc1rKQQ8fQkpfpMJmOAmYqWPmPx8ahUN4VKwmGPEvvO0
omUDirgqltdRgCx6DlUAccQ7nYHT9DTEyxYORV0S5jZ2otkgBIkhSdzEhpUlsY8oBHkdtcXELF8m
MoFQVDdXrjbdz4VFa8refOb6UZQYdyYDZtYBiVSEa92bHhmGnEsw6ff8zN+rWeCHkSYFHSgTeR6h
KzQlY7+qUY+4Vt+1xkfvoVFwhg6WLiJFRbz31+E0tJSMr7dR1mpi72qMySJJbQ2es8rU6H6oUAf4
m8H+7YnPzArFks4lKmNiSJHMSZZ4oPGzarU+lahRyehWiyUfqAaQPywe6revfk6lvn+8m0dFnlPP
8iktN7wW/72+0v+9f5+D5eKapM+F8mfBbBpM/VOrtgw8rlDZ/hDVA4i90oSB41XbilWEVgn5r/oA
EsmUwHq0mhklQ9uEf/aNF8PH4fEcSLG7dsOtyvn9BmyZp4WQS8CKGIwfb+UxllhuC+gBXidxebal
rHxJDuzQXm9twp2+HRz83a1shnKlmGywBZ16C4SwPVHwGSW/nGeLyJ/PXMFybM5koCVQ3Mf6m3Ri
XXR8hUny6dEcLVIS3q90dnTnb+YMa9D2Yl7W+mFTAoPEmYC4kadRehFEtUHRfOROPp1cObF0sdok
ysLlUyE/X7AmWjbdbk42SR5WfNp9UHMgmP3v+wMXrII0U4vXSLphl/cv5zos+u0CucJdrom64LtG
YRVSmaN/1fZPatH2HpeKBvFD4/7zga2xHW5XTGUBROWvq0BI+ubi0e6Wc/1XCUzGPko1xPikBCup
qzeQm7Q6PDCm2pQScOQN6PSCgFJ5Dnc3altTB2KOGvq/BpNi0As1P+0pz/IbJ6XR4bKy/Yxt6SaI
/+vg1nZbOF8e+3M6SDGy9sreR193BWQMoc0V8H8wd3oA/qOtxgZwCJn0UqlKqhpLhUog7ZqGRblA
396fT62i7nniDkLAOoiGfre38V/0jITegT6aSVXkQ/sGDDzys2FZpz7B/WlKl5PbAMh/3+b8eCT9
jo7jLyNNX/lbpkTptn/Nt9xOnIq6bsPdZeM5L41/2BWYJvyizN7qNSPoAaIMwl02KXnswAoPDd2c
sC2RvtXyLNoL/omzRLHyMdjIX0cGX7RCpuXkkH1fFC7v5Ia/zPAI2zBd1fj/iuuv/bxgeZkSndKB
nECqE9f50ne8xLJgrrYStS18G+mKQpou1M299C19qo1bhn/4f4OyymKPzNINJaOljegITHqETawZ
2D5dXK2w5VRG5l9dkbW5ePPNRRdUCKWvYX8LtUCt0U2IrcgKihQwdX+q4mE8Tsni+f+lkQ3eMEJh
v2fYfqHA8AYfKlP8hr8+YMbnw+ml8QhX2lwWSUwRCAk2p37E9/OsNIY/Rms5u/fjFhVzHJDPFwc1
wS2Yxit+m8bRkGydJdVZqpZLNSCgnSG2R6bhm/7zHACZZcap23TwIyPBGHB7LsJC/5ADAL2uXeQH
Q3wBGJtzf2danPSbE2wmOFiB0Rgj2ndSNH7Sqk1U6AdZ32452r4Uh0uSjrJcYgRS0gQiKUeX+Lea
SX6T593Cezz4AqMS6HivZbPpkyw5ELaGdg8jo+vPdT7g5nsHUuvYor+II776fVZDMcEOT6ocOFoW
RO+DPypCROuAsYK0uTYteo2qpCWXPzTEoZAlC0FfcwZpRNouh+iQPwKk1l/qkLiJSop3DKBZnlIi
eVRil0Ua0rcAZ4+Q/wdiIgJAnuEWGdze+1ALMsJBVj2V6BznI4wj2Bxd+NnrisRKJPEOzPZkFnyk
iT0Y0aALMxsl7tX3HUazt/49uWOfXc9xscbtIU1p80K8yUgKG+WcG8boKRbnvoc2aNSFeYhbtBkq
tl+ht8ljIAjhU065kZYds5NSaZoT+YB1aDaVKDdXERN9RNUJXRYBzgSes0EIRal9htSYls8Dpkge
4aDwtWqa2h4DHjJ7TXCDCViwkeA5MUfocQumxQer88Gko2b42fOFXb4NVw/UK2RDxS1vvmN5J6EX
XvP6hGVlwaMZft7KX9OOtQisTmRpjz24OG9IqSg0mgC/A8n67+2PYzfDs2q+ZBE7alw2f9CoaRRv
iqufGcCJbtcdt+sHZwQ3Q2M4RR/KxLuVO5dro87f9qeu8pbAncDvOjZMLCsM3hOHnoyFyiBkLNKO
7FQxNHQnqafOfVty7PCGpo9A4YG7KmyIsPe+ezh9VfNuiydaiSprGlH6Ied9GvAkGazV8zuefdJr
Uo6Lbz9wQ111FZpzNQcE+R/pn5vcE0medyfsxYkZE2yErUP8KdzupKJYNXmwU33JkYyfIwMuFjkv
cPVXeKeGHlcAl2Oent5qWHSl1xjdS3dYns394A6VDiX1flJVUxdFjzTqXExKfwm1rOYOUcU/+BL+
hM9MJwxzppt4JiMjB3CEtQ/RNI1PQuMI0B+e6cszt1s20ye7xpt1HLuDY1PjBnkvC/+ebTi2Hc57
DxFbExyDCTwNYqeHxQ22Yxmx6r4Bd0SD0iSdr4X2OC1dTm+RqMW/4RE9WHPjrkC5NDcmc8wgZBX6
nDukYvmtAMPromyKrY7pEWvq1e7EsY0t0pT2jsu1ikjnz1UHu6Cq7mKkjL4/9wXJ8DPC4FpppM90
y03CM8IkJanlfI78osD0q5sP0qFjtFr2SWXNuh8O9TAAxF+UoT1UsHnB6CfCsMPjwMZOMBrXVurE
kjrEtrqX+W36GfVVFuuiQQ8VCwACZfmTEpNzjHDBGEvNPvwHOyyBsvrJK5uE9tMgTWtGQJISTypv
6tTFpfSKhsGjGXy/IAk+6W+GVR0ydkaCA/eLgA3mD/mQr+ANxndlG4IxLBy1kuDlGuEkxIA6OVpw
ksy2bQkd9mf8rI93WwToEgmmKVSUzrBBkkhr/jr6C4/aq6p53fJOMzu+aR9YmWYmCUL/7wtJiQU1
kjXLYG1qSmUAwV4HbYM6ed1zSFH/LJQsWdYTkuzR2iWz5ZWlWia/vVs+5ZEIvRBjA/0K7CS8NwDr
8BHfAVY9zrJWrMVlZWLJziLONbUIV+xwnRqZm7+FA2hqo4EepTXlBj0WjG4Vfqm3ZTGWGFcyXhbf
akA9/1KOVGkFbz8TmvqdmUmuvg+fLZxtrkYvKIRYgPtdGNtaZKBMcCrRxu2z/KJ/kQ/xY9FgPEsw
tacuiAd3aeOSdmrn0/7RsEqemKC/0/um0EcC5A7j04/GNvEEl7Yulb1d5A6cfoJ8SzYURi9flADm
iQiTGjbVOxYx5eFFJ20h/WQrJ0JeLDxzM3fp/aceEKZPvLaI1Tp89xG51/NinEGVaLQA2XFV6M1w
QzG11GgrhTdLksp9PMzqDkbZ3D+PNh+2qmJsnD1npzvpYwI4UF9tl19Y/x4Zte6Z7q7CzlTiG5BR
iq/LmDkpUmOST0WgJ1eXLg/rKS2kdCQWbNw2XhMx2/osD2+kyPrfVnT7ozoIH1fwanAyKB597Hhk
MFW1KPU9Ooh8CW6p2pMnmg//2AUwU0g8FNRTKv8hKXlrElYmgRhMdwdzyhbsPL8p41N1yIvqn9k/
d3j5YDlW6v3WHLfYehrjHtLMOfPfI64/usEIe5BMnRT5nOjwOAWuLSg+nClH5FqWeZXektJrC4N3
Kq7nmodpH9Eau/AWix9QQJoTkofm1B6WeM/pIHtdw7F3OeMhLohOcgRS2/r/vOGScDLCGmkN9di3
CVwXHcerlTBZp3BzQaYWOMgkXmoAnKg9MkZQM8zGcEwvNCS5cGfltz8lCdJKXGgUGzPP0gvMaYmd
fGKEHGlc5zyShzW+YoLmKBPsHd1uNmyNj7y+XPfe9y1KNiH1UBZNhPKcywKleGf5O99lLk+rrX2p
LkDZMtTS2GiZ0Ig+vfT3osDDRBiDQ6cFJxIurUp9XXICubLU+z4gEeUtHRW1QhcHlpWVE7jkJSO6
VPu2NI3506HvPGtTNgtw3IWIFvO+KZTmknHOwTQAfdXYaZzX/KFauSNf62xy0D+kWBEOHVPvVLn5
6jAXkOEcnvibdvwgpH53nXq0MhuiywjzrLz18nyKRMjLUD1v201tAPPRynCgKvNoGKdbM0T8QlZ+
1NdcNGzSiXDvBaY/DCKn8eMI2iQxsXem7JO1YUNEUTc16JWCR/r0VWS0jYJhu2WX977K0NtBfttA
cjz1qXtMVnlM/dJ1CYtJPePzRKh5o2MM0x68Hygm5D6L6+7oyPPHx5G4MEQHUw0VTPR16D8ca6Wi
D1JkyY8EyNa+IA151/PYQ49s+Gzs5aFjJvpgtdmzjAVNcRtSDa5HFHz0/ZRGoCpv0B1fryh7PUd7
rYG/FXr+TUjJrMd5FBt1nUOVCY8dgQW+9SHA9T63QPEa6viQeT97Bo2YlwqOvhZH6sWRWm4Cn9Wj
KyeaQ78IlZaZORIm+lMrih9Zoj5TC6A0lDpHJWfQI9Ubgj5HvfnvOQLCxl5Lwv/r+0WPoHR2h/wK
JxLdPfA9QLWKuMqBUxfXPkdc7Q8XZ/zTcF67iwFQXX1uByb2QSSp7T1ch9axWH3gB6L7Me2Tqyya
Qc4CXoGAS2w2e75hflELZbv1zhi644J8xP2/tsP6Qu3+Tna24xdu+MbxSVQwyQAJJJyKaPSmeHqy
sH6ythkTRl1zqEQV/GSKofRQaMu1X09I8kfXkPIJ9/RvDnwHKDV5NWQ8UWHv42lLMtLyJa5uEOvQ
A1x7loB8eE79laMWpVL534GaR/bGGxHkhuxgsaVpmbNk9WgfAPlsHdSIsXgqOwA7U0HfL5rv+1jB
t7F7f7dXV4MHPK7or8TUCygih6cZ9pnWYfTTfO1yFYalyGVd4ou88Iif/ppBtDqJgdIzvASqRyux
Gf0+/FcERbI+QNu9T4+049yBxpCgF55//BHbFmHJVSOpDfTGCcm/GEUS3S7nzNKgj+qGJzVop2QS
VSgQ/J5HYFiP1iLd9fBfMK7zW9FaArUMTeXSRyvSosOccgrYZfd8edsWVarEH1XqyI5PlbBomqBr
k1Y5GC2erpGEQ8Fqz8hUEG2qaYOnUh0jLeKKJvJzLcj8ox2DXJ3RB5y8w1K6mfO97MS5U7rTGG0z
XeExb5tk/weZSYioBXNN9wX4dzM1gX9Xc6buaCXbzzFeaH2VpMTcqU5x/nXWv+PDe1pYItzk9BYZ
3x4ZB3/mrkZdYQcJK8NbICMCSc6nXNXbWpPEvGXVq38RK38BtZhSb/u8Sp2bND7Z5cjrr/kitbHl
eCOAGcbhN7joeYN6t/jEKlF1Dv3xXm7eEtMwOhnZlW9uypEfNjH2s9ErrLerAURGto0ni9G8L782
NzK5jq03b9QK11+SKUVQgAaRUc/vOFhLx5RQGdJmm2LCKV2ozTzp80fRGtJh8RqGu4IzDDljOZpe
RYdnOcAEZv7JkkrOWoABYcXrMFfBWbqaIqflUPPlcHkEgkIjmsnlnSKTPLU8VvFw+eoJHQjtnKTc
XW58J5pyocRZvIdw57oTAsd3wqsNXat0M1EEmNxal1z5jfnIMK9bRcJ9XZIxV6S3ljGofHr9Tapo
5HBckCPhsW5vRgAuuXu/3JJp8INp7txDGi9qE9IfMdEvlpRRxp4lL7hyUyrrJpePyy+S7aLd1DJx
6wW/kq938I7CkQSRaK/CQGKxbwAFGU3RVNCAwJYcyLioCVaczx/rpM1ylCc7DrnD+B+LhKVLs0nN
lLbWvdgaoJ4BSKFmhdwBRdA6isP7mogamDxKlXVRs/kDreNkRYlG8kv6+8Vfugqfgr9QrzJozjg2
HOHehr6plwe8PUwF4ZQcTuCz6vUzhOduHgorOtzGWVx+bJqPSeesPGtRkQ9/TUTTvWl0eee53bwf
cAy7i73j80EaHj0Jj4x6vX0qJLg1EgJgfn/1uDVfeGpGU1vbuTFKykqlhXHrESY7TGx7Bt9IhnYi
cWI8iQXDhypPA4L9nxaDiMRrYy8eUJHhNut9oDICvAE0NouO9L3a/8ViyAOxcI3uf2npOR0AG3me
RwyBfLe3uOsdCQiGQAQ9U59v7z3Frvus6laHNyNUnNKk9dBUgDuq17FaSm6crdQjIkETbG2iIPq1
T3hDKuR/sp8djm3AdslMThVSfw3Nvj2uNMAq8hRnD7FsDvgf0nGnSPJbvBv3wjho6x22gp6hCYts
XrHLcGfXXhqYD0wvmRANar+/AUP8hp92cWi0AIpw7w0250YsSvgNmIT8iwyPgSLjRWmFQ+yTE9UK
zr5LI3iRR0GNqATGI4p2XcgqD6izUL9hPSPpBD3WF1e7VWy+XvxjBGSaA5ZlJIXCV9hy1LXjyGuS
xe5iTL9W9by6dQWb72Sn15OgGjUcR6/HdoAvtXUhV20jDq/SWfUJNkXXvG3XNtO0wG2tt6Dkiu3i
Gn8Cctp5sQLysjFMSzThat+E83Qa/keA789jq3B6RwGKVaB77B2zN2esOBpox1rMe/rlSna3NdB5
8UIH18Aj6l/daiLoTaC2KwyCneNRVFZQroyyZC4tI3OF0oJrNjgyA9xAzJdJ47BAcKPhcbSGwaXm
0gu9aE4kHJywbLLxsdxqU6AAM2oMg3s3zFdXPRMkUh99OAATiqxSY9T2g3UgiB2O3Bb74Y8ON6/x
W2714Zn9XlXsERXzyI8g0u6a/dgAq1JDhxfDC7e3Me5f9JuZQ64/PSnud9xuach3sJO995UdIabX
ws/o7KjQCfSWvJIc04O1pPfNszCeQMdDo2vak0CQqwHG72/ZjVtRTjaOs6hQWdoErBN5PTOEY+0Y
W6YiVeY1/7YJwFokXNXKtUedyiZ07zF88CbSC1W2pbFFUza5xN7Rh3iRsk7lfGsEpFoTRMyePV/r
PcR90TcmSU1F0MxjqWQlhJpD7dYmqRFBZ2+2lMP2AFGNRVOmj6xvlyHfM/cqiP5FvKlBnQAjL1Ks
uVKTVCxd9y29GDT4QmfRoRD0WmGzTxSTHrpaoyN4/qLnWUuVwnLwzJmCGuPVnJ3gnhLVqCiAVN5d
4OBOvqVNbQPNDVJNV2w7lZXGuJSRe5oWnTw7rKIaRhbJ1E1uuRptmtoRiz4XopLC9ykWVpPf2c5q
lEqOf7OCnZv877Ys4C4pVHSc4MH3HNOQP+Tj/sbMfyVeppLTuZFpCFDL7oPAI7zWx55h9ZqPjz09
Iu0yAxKboGFkBMdJSIjJpeWWiM3eT4oWhrfEjeydhqJSH6UdxvPnuvuY94xlAk2ZjTrh0HeFGpjd
oihFF+8IS8clcsFiAgLbSfaugPif8Zmkmr78DB6zY4iG1Wh8r6H2PA0Nx16nJuWE6VqbOFGdHNSx
bS+Rw3B+rr/XHNk7+Aq8qRqPuGh0mVMzILXTHaBXkL3L6imuGUw2qH7tnars26CpGyadwnjPB2kM
dpgGlYHt47zySHKMefj2rkW8bl1lS/gUcHVlfpm2P/+X+EnjnOwj4iVPUEFOAfuF7vpqadQWkICV
z5DwoTEwq5zpy1Npem1lZvW/FwbF9kGOifTVBJfLWavsp7RB1tWgNhZnlCktJE2CGgrOrFbbFBTB
X10qy/fgrSh+iPuN1cV5OoQjp6tKOLmSrrEZIBfIoeRBONRdKhArS5CVnAol+1flvGvP3+vge3+Y
yMHyi4UUMbGhg8ur9r/q7ofu/vSnH9qXMIC+GNvKDuAHrr4xH4+Zylagbh20bnqr5IYxDRflfJcq
XzLku0X5IaRhfIM0b8j6k2gLYbg0InQXaxe+ReY0gkTXI/HFi1USVcFY5oJP7Nstze3M8SxfQOR5
2X6fXCt9GsXTEvo3st6jl0N37OlYQIPR/IFNh0EUsZaQ6cD033IhEjoSVM8khlAbOfBiNWJoJouW
cDYRnCUQ+QPIiQB0Zii/VPGBfmGG0XLVmsUG+ZTY4L03v+A0paAVGxS4S32RL+PQS0X5Gm0Kjj4f
i+zNYHcWHnXF2KQoyKBKOiWRFpjXB60qnmRJbNweabGi8a64eHHRvwzBAELTyFiXWaEK0EANGiQB
E1DeahfTs/IzThY0eWFZDnh8CzMsGC2nzWoYl7AU56q+4zIHpuCwfnulORDVkn2bFVzpZFyNRDPf
95l42kfilhjlYMN+0N1LVDT3VlUQwQ7Tm8+b319853Y9KEH6Dcp2wdxP+EYksHd848gmn1qgEmBk
1jn2D89mvxY/AdVHfpKAI70X7h/U5tC5V5jl7SSArlt9QE1y6fJ6MOmR7CBwaGQfoDLkjiwKTWXT
YcS7mBrOIUtLvAhfwqlfEwJ6SIM6WAlXuwxl+VUqwKvLmx/u5E9Ftgz9FNcKXnt3+nopQ7I8vemP
xKIN7zzEpWC2PWYn0To3ZFUrXeEwh/WBc4K9J+q0Q0vRsOJ8HQ8OvztsFNlpeUYhbjKLC4V5Hr10
opzdv6KbUtuG24dLEOwiUXrBJhHbdVOIZVNtqJmEpDxtMR2dC4oxf4gEhN6GbGomBNEXxLRSMa6n
FKfavhRMhQOuA5t/GWmD5ERPpYYgZZ2CmulLp4DMhEQxK8CsorYpjRDB4xogmjFTjkwLBFOSGrA6
lbTfVCVlJWaTU2gSexNxf4UUgOHZl7T0kx+IXu4o3CJndwk7U0MIUBILLtyTrIjntoXFvSF20Kmw
fcqJJiq2QN9Nl3CCecgCMtQNVgnJKXffraT8wlNv/QDqNTFjgaUrvu3fwPrB/ywwJU8X/4LlsN4k
cXuN/+Iy5M+THRUzCzIbDhBvKXnfTJs9P2RrYKTbwRMD4clDBtPqHhdjYd2+SBq6+nMUW4SnCjje
/JckZ5gqFfov6IhO3wRpWEi2k2NEfoTMg68RRnQ0MafpOj5OAM4L8QehgO2JjLwydb2MK47v8hgC
EChXycBLLVe9SBnP2NCGD47Xk6UKJsvaP9ONlzGBn3OkN/DNqpbYtEcse+g+Q/eVo+p5xUbvponF
dOB14/BYQeox6tqHMiRw0fUj39/hlqx4wx2eFt61XrrNlKtJWi4iF0ZOTZ0o7E5PIPAFadFUita/
UOnuaqP4e1XzpJ35rjpAZhlMGMWk9MkaRgddIV4KNjdhAJ2ageJRi7QPhHIoHLfppJfmvFkS0U6L
Af3CtdE7eRalPLfp82VLDtX5ErxztZHU8zZgnNia+/Rt+LOYO394d6+Loxx+7vl+E/bLbBSYAB1o
uBjizXG3fU1fNEY2hUViE0aWfM/QRPkHtjHPalHQ5SpI/exAXgfn7Lmc+7i8d25zF3qrRYAzuWlj
DOaI2esf+6M3iQD8daV3CDEz51CjLsWOIfOGzw6ozSalozpkTnEtr+ln5XjtUJ3JwOhoNGKZLsNT
Dau4d2TyCQ/1UqIPO0a628q4Sp5cNwLeJywsOfN0/jW7pVIMoHRxofxvtGHXFuidjJCIk3vWUCOA
quwWWYn9LNb+stM2fkEreX+QxCz9710SowYkgnzwcCSFsN4Ooi/IWlCv3JAhfXh+TaVjHsxnOaA2
GeD4M+AuZT3d/TWkdusPSyG/s5+dJKRl22mOf44xilngR/IS1MfYgp4MXz9fOVR38DSZ6d4DQ+kk
GUD1sAP0+xfOKRJ8ikV8haLpupY/OASf080qhVqfUlY81VWM9+wMaiv2Afp8oTqvF3pAa6cU/TbN
GNh7bPuljh66OUOi3ReJ2twFH/XJuu3LZLh4ck33m0zKxT7uLP2cNWM/SdhW3gJgVQ0T35Y57Jta
VxcYJZ7+9c54KLfbbH263CoRnqcOY4oQHjPLIXN/fg9uOXM89Q9kR2RoOvrHbIjuJEzSB7uz2KeT
2bVifOYLwuK6klwb4HqHqONqASfXXHcCTFTM72b0uvcj5P6pje/YA/gNJyZTmOGx72fcAj5t1mN/
HTHq3XqsyyANlrPLBZDOXrMdH/MPqdFUPjwjP8NkZ5ieT3mzq2qRNLxwPYK3hD/JEma+Qmdtigrm
tFgJW/SXXKxTYuy1RHm+4hZb0/vREREP7XijjFCcLxT2V25zdz1oFRitRFPl3IPpYr8+shMN9F6Q
IUT3MUqWxMe1OXtxW0vVM9oF0HnyBibMqeupJUqh8Rz6PseXym8ZjYjHQ8WKOobVYVlz/MMalR5i
l0s2gtiOjaFef+ntP+8OQj/suWqgiIy+uiv3Uj3TT06njXvdoxSdKjDyhFkQg2elynT9G1BEgQzo
Xv96S1UXU1/WwnsaVkg2b0NfFyNplGK0VigWeuONa6O156Nwq/waQp49vlIQDT6dAl1IoNSvJFfD
Upg/dceTsuP8Tc/CqpP8gvYu1T4VPWpL9qUxw25Sq1PwGabr8gobomIt5qw+lEZf2OtJsjLpFGgG
whxex7AUMkLl18+TuRR9xgFjd076jPf3PUKWdkUSuqmN/M1ExfxBlBpwR4qqMExyIFqw/hu7WFHu
OkaLDdPvtUt+pXMkwGq3XgdtklBRiA/Of1ZIKtgdOnzoU3ouqDT9n2N2esfBUYbQmtd0Nd8PzS/y
NBE6GwVymyY+3nely16FVT1h1hu/hZAGF7NAY8sWzyF2LJXvGyb/ilRorkrqZwSEzfdqPcOQpvwX
pv9pIkmBItFcWpkYBvz72Qxk9Lk0ilh0q4TIxFabMV0Pke2Mr0vnBDmMutmW4q8oIy9lJ0bg4h9Z
36g7/Phw1PwjJLFRYNJeFVar9y7Psb278AOAsosIMClYsSgPFfTuenlHZNMPRggdFHOJ8aFkyOMm
Y0TypGSjDKU437Jf4rT51lj+zcEI67lHVXuqkcT/z8bVfMqoj06s5TA7aP9gKENr0ry0maBqPK6N
BST2JIdi9m4cVXxOn+r8geeOIhFIfHmA6vXCfoh/qzgd5Y4QUNlfrpYlUUqnP8rUA9UEZATHYDpl
HN0YVR4iJOFZ59z6kyzi2GVHzUH6ABVuR09NzMeZXqWL/w1R7gEfsCGwhYRvbfp1eRvmOduobtqp
hbVdjelR+Q+3BYDsrC/oDSNzBxQZHtkbGc6659PJw8PcJ0cS7twafe3D+20SWJYExQbvSlG+346b
J10wk+cL/YKSl1YK4e3878tnkdH6xetjafngiOk/nVrNV1w46lI6QWpe+u8KHNV8nPHlVOrALaUK
eN8mzkQLw/ZX19qSFaZ1ao9fuDBd6z7YPN3EGQAFr91eUdKMtrE6WRcI18LEPmcVXXawrA3Y3XBm
jqPN7Dm66P6b7xCU7EMNLGwgBID75EPWtDBZqCt0Qs9bASQeIVDBc5zMHZ32MYDirLhzMhIdcKEi
WLeFrviqi1VdG/qtJ3QHKiCr2pAZL76ll2wFGLaahJk/CISMzTsowCiXSQQjD0wD8dbdFs+66mvq
8PtYRYaEiGqkWViGUGeBhf3fDt5EF4f8Owoqal3xQOsZxKUtF8NcgLFeUYpHhtz60P/a7Zy1UYNo
ruDxQazVkkyxjidEA+J8Sb7DK2m718Z1kitaAQAqvpdoe9L2VKwdIpmYjXAyUCyoNxiitOpZEkaM
1tM4bzxnATGRqWB2JiKX57Hz4irMM6uwAegtabz2nKXOm3q/jHrWQh2KmXa/wXW9jOQLjIMn1ISN
midpqVbfN1m45Etq2kXNZG0/R6DG2SuTJ2Pum9bQE/2i3/uqR3nPxOOF3F7WKiBlnYJjYgB5I7Jo
GnGOzYHjl43IvxK3bk95iDUgUbAaty3xl9xL4C3qrnmS6OgVce3J8NKc3L5yvAyO/7FlOMr0+mpF
K8C0zB6tGh5MN4pT4Ve90HKWUjaRq5iP2zyiXNj0GnGiAjdALh3Namzn9RD1ZjmYM1EwRysrldFe
vtGRGRJwJFNTCgRO6D67b0WP8IlyHDcLxaj9QYthjZKiS6Hf0JBnOli7sYo3E3TVmJFqslZ6zlme
yuIM4ldB1aKUQKOVZSB+AJutM3qGinFeuqAgm/+oFrqyWnjM5tyl8J4cKY3FFjbGgHLRmxIT2d06
FEn9EoAa1ItXvJ0syl1xRcVPbsS2+y3yujT2lDKJ2pAxuGIXe21qa8GZXZgITFUakAYPC1jNPraI
6h598P3aRgvsPDXub2Al8iKnZAZZQo/CmhQ1Yf8HP8VQm/90nbNxhMJkju+J8FD5zoxvVMogHy6h
mjkGzbFLBRma3baDjja4W0OErLT9YO+QcKXFboFQmmZQWJO09MyUNMWMfALG8gfjKe5zLrCx5RHh
J/LygWnE+gbXzzMDbfAimdJ6DaqoreG/hJlhS4a04ZGENw54QdPkLcX2uIYwZzuV8nkjiRnbPmni
W8LfVO2+df4BJVCLA2CnfgMDoNhYGPZnYWSogev16IQSibwlLwQz6R6b39le1DsFZqg+oDPwqYjW
HxmW8e9NaOxpUaI6qeYTNDeRv+n3S4wOpeLxw/MHdZ53NrZtFuCCwDOVXmzMc+pv2y0bhOPFYzcP
sJF8UWMHOtTZE4Lzp2/CM5Pz7gclE9WNkPm7wl6XObErxwAsgKgvH9UxP3r/sPktQVdzvvRuT+qL
iHaJXk5C+Z2dZhAYN9ujoFuN8q7AcFmLSJpBZ+MeMI6lDOYY87mqA0dDj00xBY3R7wvOlRnBWdF9
5dr7hHfw7b2Le2T7y+6K/0Y6Z6VR70Ov0ku7/lZeSxLN3za0COBlCr5xRASr+2YfYfeZjQlE9cbT
5Pd4iuJ0eMf2paC8Peqsq690bVYr/Mjb1fjxz6IxWyou54rGDYd2be+vifvzZiADGu80TtCKzuY9
IrsrPACuHKcxknnnvnQD9PPt0qdUQzAQO/SY3O3i1U+hotbvLfS0+9jNHQIWsAg6eroBpJMrfMg2
K0ke8X7ojJr2gungl5KjS/n3pocJPlUIcoABXQzZpvc/Gb+OthW5Ls6+yhahRuSQnKWwTjNxkr2J
cdotYE4zukboZDKblquClVcNYzAGLT8iCw1+O2MiP3QJwyJSoUZs5woSJ1wuNNSRqWD8EEqtzFa5
RFt0yRDyJ8z4mYDm1F9C0R56x1eygXCuHbDpyhs6Ag/keMel1cVsp3Yl5ASXs6FwWu3w/Sypho4F
q0UbxlqtdEODFx03AJInD1uRijZcZKJetBFvQffrj2SBHWeBb5j/ychnGWYmprGEwBniZZ0jiinn
H7aGBnZ6/NCUfGatUAOaYep+jEIrC0XNrXYX85MClyO/bKKBlUeDalxfS1YXxqL1RKfYt/j/xE9R
P1HqtHtkjPbnJIOP1FV4TKRYkBaoTzZgW9VWzb1GMyE54ddpt7e1OPc9y+j0ixdvIRQHtEUgHs+u
343ioGzqrN6bd3yKPq9kWSxE5jA/7BuyfltMDIGyIuaApIhYXyKAGIa31EiMorRl6tMWwW0GAKUf
1ObJerZWMvRGfY+R0J//x41ncGSNMryRpTmPzyK9M3bt5aWqTFjTgb+9xXIwurwBfa/AghFro9vn
hvw0IGVxKTgQISujz7rkCzZZ07bF+ZhoNBf5P+H8+7j0g0XgvRnGuOVGgd2t/vRM+VLGEuudTUO1
6sFuNosd72PIH1nptM302XolEV+3Htbi20WnYBb6JgXpCAyh8da5/KaIJ3QAoRKf6iXf21qWQRJH
2UJRAZnVH2p3AFiNp8DJ3cNy0SS+punQc90MEdJwde0QgYtvtnuCWKMK6bYW7vcvID3nkva47iD3
GEhaXI5cyMebY1Oqzgqk8SWCLABAu34UJbi+P9Rv6BHC07O20wrQx8tszDNOeU8+oZeWLeaUCTTj
sXlK7px1Ny90v9b7UqqxVpsk/Pl05dv6iN7D7itC5++xRVakBpKZQ4JlE4TrBUpdyO9z1qgmsIvU
gq0V2OMBEXMDetb40nIVJ4iQkBFYoOmL9nwHjEPNeYaegTZIXhdysr7cyXzxvHHfniHb6+wtkygu
mwJKk5GioqbeHUvbSzEOmOKd7Ee5WNeTzmoWtVkhxBikHfWO5wRBh2j1CjBHwWcaPR2DbUX1evv5
sdssiKT0xT2R/H08WZ83Xj6rhX7SW8nVMcbnnbo4GcEKYFDrjZ1GFIq9SjNIbmafGv85oqoXtVwp
l6NezjwTxSU7l3FRdDyP1SJyBLY6hBXgWH/rAH5wxtxSEUvirhmH+XXYDfCv95IJrCNIN0e9pUMq
8Ajfuk0CTbVuzi+xExoaPbmJZ39UWCQbaE9QnQtx8jYOTInwK2eLrxjF0O/Y8RwreOsCd8bUg2jP
9g3pBdpisXj+uif7Y2k2G/UhHoXu0U2Bb22zlJml9jZrqYdXMxu9Dat7KbkcymvTB4D9FTISUt6g
mh18w+kSGI+H0+RolMx2pfFWptjrznKajHBp9uPv+IZkJECWyOq1MToLZmuo5lsTeHxJcuur1COU
ji8gQh4KznsgOixGtuk5DUoxhaOHB+jULQdmXOkBwStVMaPWXmCFb/aAl1yjdrpHlTBj+OUD1vqn
B093aKXixRWVI6HHytVl5kgJ/VW3BiZmQED1tgZvIVJhC6g9Lv4NUF6+3txJsJzboYylfCAYSrRI
Y6Th86+HH8OQISheIwMuamG28fx4vUi148pNly15237/AVbfO7gsWX7xUozqLyzhgqUqicurFzGo
rMslhX71Vz/qKGPR3RlkuERdcgMYOPEj8W/FlwNyqx+WGsgkRCBIHVSu3VmsdiBkvaBdk5+kRpAD
+fO4Yfv/G0NRQSXVg6ezTKuJT+b323S0pY0gzocXxTj8FdJId86rnpaDBwvNhVx/3xvo+bdrzHdp
vO3loRupENA9sEs7OVEGoGqlxJHeiS6j2IvcYlfTZuSiAlQPugf2LVB+2aArTmCsV+gbfS2JhfHj
+GeOmNRKldnlGach7f456dOw4NyGCgFAzmw6MgSxKtuh3x7CBlbuKwrxgUAWDnbETNlbqUNACsWs
QBIq9glOZl+Ab146CvSdiTWReUv/lg2Hv3RmZUiioy/9VvByu6/C5CpAUwOWHWP53xu9jR/czRpc
nbHjAUL9zbaKBDV4ZKxuxnxFZQUnK7k7q5Owg5A6Q220CSdtR3gjTIkynNkk5cXShGNfDjWcxltM
GBzzGmkz2n0xtGTlRVgrl7R8ToNPmLEhSBJqD+s8vYHIcxc6IbVXtW4xTGFDKnT8GXdxrz90SqAn
6sCseK07jZ9VUrD7STiHQZl1zbc8ON4LSZ2LULDJ67REZ5G1pC/pa/QUacfsA1zilPTFOXAbS7Oo
w0bHLW7nVmcSM0hZXvScD20RXzEMO5xoQQwRpv83znqmomO/ugii6Q/HOWGZSK5vaNMNUicbIPgB
F5HtoTGBBljdBoW9r4tgPSTNajuXVVOMjOoeY3jeCFuqn+2RQn79gNziIE/V2iCUjF/lyLSGjpGK
9vfOPDixwfge47pqw2dQo/Qd42WIPxCnrZlpG8hz2c4pkxfya9uwrQzSrsrlzzNAP86OPv4LF7Bf
gG5aj5n6ReV1+d+axdYTWkyPRo0vPWrgQ7uSeNOJkuMAyNh8Oeuso4dPFafMa0sdy3qotNAiYMtR
CuKXtt1SyBVNzmErh6FBJQCrLQCpTbTbAL2kFZTNTzBTmqMEuOmJh9c2XXMg/SSl5zqcUwelCu+x
mvQNn7imQp0dwsGzvR1XLrKlRFFosrxcmp3mgWYKl9EiG1Vh5eA0hvcwtHor/KGS+effFimz4Swo
SnndYl+gPplFBlcRLbcy9hancuyaRea7SHaJKsf6fdYKkeL5PYxW8HrK4IptiVn34VItq1hQmueQ
SOKe8xe4dTcFUD1xMqZySXdhSDYg8jty7X2LzOm9lSs1QC+RaKnSgiscLEXlTJcdOlLZbKuPIdzt
rbyw2V3PuQ2l+WWiUqEN3vU2iYuspidIVNav7FThy4utAyiROunNpqpab+EV5Wbs880w70/eLSgo
UzNb7h0Ql6Dt11XSaoGfXDe7b6WZ8svoLRCrE6GrpQsj9ImVAhtlHXFlRlcuipSTNSvgP7ifl9rp
OtHRHBDwt74bOwormsXBOEi7L4Q05zMW3IOtxq4TTnkkqHh1eMgFHj1Oa2hj1eza2T9qqHa5afPT
VAmHpRDZ9FFB99M5ZSSJVLtzVr7kk2/Za2Teu0tKbSG2KfQ/Ol0xBzNBKvgnHhAEt10ptbM91EVR
+d8ZmKXZRjLh9KyTPXI2ZREwn6imGEGo5N8mgsGG9g4q2MQXsWKLDevuHmu4sHhruDAk0FfS3/HF
trL9wyxqYWtLQPIflQNS3HOjA/2SsLAR7HLG9z9RLA9l2UWspoM9KZSZZvWV4p68ASsu0Eeo4c3d
jBteJiogPyDDqZj5/zecBJPjnub/YlFSIt6bBZnldCqLjQUASN8xlzGTaJZYTSpyhkZ4b4cDE2Dd
T+q/E041MAfUnseHff44gn+3gVDo5IMskrNEm1U8BcgU7Y+Hmr96RrtzWpeLzsHL4LtQyuHnudRt
6Y+ESaUCaG98Ef28/663RZRFgS5YxoJgIFAlSwqVKsyVeDviBxS64kYp+pwvzhYShRyctOuIL0Zl
gjZizJbKI4LYJxTTj19GZ8K3HbLLHYiXp4vS9TllU6VUtMyO0faq6gVvAy+nUucXUTgiVj/n0Oh2
XTkQfW0myMme+JDSO5LvH6IPu8db58/Zi8oCg+hFpkdAIwBjPz0+QM6Yw5n0gK42mQboM2tc+2Zz
vce2oNKaRlDslDn5kQ6vWjH+ZyGg1gqjZnBO/JYo8y8OikKVbb4yhPzh8OiafyXsQO5v4s9IoJQ1
sw/8+uve91Onml7QSkg0JVaedF4k1J/ZZSiJMri1AwG1is3J2egwcqFHiZhJ/jQDUiGGgXPHQ9pA
zdehNypS+EWzviXHGJTUYUyzSxF9D62mNxPDkwFgsrAF8Niqxu3lX1vFeP6Qj4m9nnUxPmIMd4ua
QYt39xeruz55sjO61vRACcxbu3wGjzwBkwgkzJjmaxYjBNTrNfBTeE39wdqTKv4RsSGK5r8FoIaA
JlWWNDV64ix+3z3vSEbu4wdAGWB501sW5hmajMVpG9Zq/bbgwwqaj9NuhxaJlaLXq7mtVnIrMpje
Rw6TL+iHpUUi51vdMq7MWSBguw/OYxHFX+nKfIQLblJWY0j9E2kcC147hV77nPf5gl8XHI7k3bRf
17wL7qf+q0ITvMyPsgWVyG3ukboqY8ARbQ4MWQQfoEBBZZKFMlWiC8zIeyH+ANcz6ycjbo24ieMv
16sHglW9RDvjqcMTDjF5PA8HR4WWJ6cYMmqZ81ucEjlffJw3MQzzNTaakvkyyg6GE1rmHbBZ7P4g
tEYrdxCTAhvytHnBFa2jDswM51H2hE/G73kiFz2tgDsCinB/D6R4f622N/R/4MddYV01D4lYi6Ft
BSBBBJrtTxW2T1mFVUKaychpd6mBCFw9tH5E3BnXp29YFFlFoZp/q9T3NtAQRC5WIxsOYxMoHjfw
lrBeFi5HYL9koG8bEr0ji1WLIOh9feJta5mKzCZ/06aOQ3UyS58nhN6dQ2Twvlh4+KYHuUCo5A60
T9O88+Jyoihaf96dtWB7qjWaPUNYUk8dAnLJBvGxASpLSn0Gy/4GeCrquU/CT+s0oKY1ljW0hL6y
UpiSKmx5ygLUiZ/BxUckGb7BqEY81qChh1zQA8rwYOAbKWsTPGUFp84XsO5TuV7L5VLDJLM2jQeQ
k72SLHOqYCyNpRtzCk5ILeKJ11gRkS/zwXjjVB1oIJzM5yHm0QMUC5bYicfkQcBWTLXQHzH/P+HY
Cag5GzsAEaZVYRYzhBVMm5EYmHlnAggT2j1VYIwE9HlQIPW4SUrpGDuHISK6aTOF1zrG/l00hTqD
FSXB7CYbIR3BxYsotkO7sbbNgsJX4PbUZ4EkL4/gjQNRIEVmg1se7gjsIAtj52HlV3PG7RWI3NX8
LMDK+YHUfTqOb62GaRBzHBaGkvdzGTEhJlW3Nz3ArGbW17ONAGnYNXNX5WoZ2BqEzeYmnpgsePpl
ocXpY0mEtkHFMrmw78FXMDjswBZhr2srWn3POybuH3M3HzjYL4vKEmyLOJoVCG8FIzVr5WKaGsWC
kKd/rkove3LosMoMe955axcnx+RY/4g/jM3uD+WDk4os1aVRcpUH8huwQgb12PWG7qFne4h39qUG
QucscIhxZmnPFxlUW1SHgTgeEZuTDK9pgxr5PNKTjwbM5UBx5klJ4OQrygD4zvcZVR0s1oQLuHyh
pkcOtmKfR3C6hMgH+K3koWV9DcOD/pZdUZvjmZhkQ+6AV/qYGiYsh+4suat8AHqFizNM3FWo0/6O
xPPzlUelbepncSBkuMS52Ct8nf8dDxz+i2kRzsdP9Vb/zArU/03z1UPvlggamR0LrW0kTmZXbXAn
OajuK7N7ZL4X+nqk8my8PL2MN2xLCWLMiGFPnJPBMOxQNpmhlsdtCJeOEKmvg69UoYRJ2Uiq86Ve
51IDPRj7Kj2k9YhCf89z5I04dJ7QsYrDSshzcrFMHml6XEngoEZ7lFjPqJSCg5IQwwOyo0DBpgCF
W6F5xk+HR9KRc1lCMbTXt2uEZ8acKXirkJw1heS41saNCBtQbwmcFZrZU4FH9Ek8mvjz8QPgdJQz
/ydjBB4cOZKIAlzDlx3GODdjW8WYilR9pW7S6YFzU9BwvCcmkkPcI8a9xdaq4t4TB6POxAatdPtN
2zoysqWsiVPL+JziGRE2iUg5zdG0jbszFnPczFhsi8cqfY65NwbycxDyE/osLZLw8LxsvvnXmnGf
gs8rDh1Plq8oxiX2ca210w2+tsFP8lcD8MO68MzJTLIdAHrdhsBNWTxirsOXmYnJ/Jy7FaEWRlDf
RFupVi+iAnU/XZHxOMfFVJ1uzrPNfI3Ah7/y6P7uOC0XbWIZ7ysPl3ySMFIKTCismpCHttDhrh1E
rqQ0K2S2s3wL0zeIf/EbD3NpHEzR+AVq0XR/83T6h1iSC6wWaWyVKY//+v/tcvldHj79Tn2S2DVC
NfVHqucY5+Qr3WKPF+QDLd0ElApiw9NTwVdGZddrjA3T0HM5V2shDUuBNxih7Y3zTDapTOfRIulC
ImVHHL7XBD7KIpY5QpZ5qWtUoDSZmSqAGCsdQKX6lXUoZQu0ZU3Lh+4EGjN3cAI5yW8IPhdsXs33
J1vrGAiQ1Lli/83rlyw0BODk5xaEufYhTDx1IdxFnJQKavtxo/kIol2nLzDiCe1N/2+Jgx+wwXuo
/f1xYcScIdDpQj3m9oikrPpiCdtWvG3T6pa9Z9VhpqwCEqnQsHo+9tfWuWODyU0LJZTEoXIsoVOD
9OTZujHp/urgPdDe05dKo6jZFx4ruAGoOcxnySb1f88WAevLLxRtn8unpir2D6jl/iN0frWDlxRY
eMMiGPlw7YPnVLuOCvI+QAWsoN+E2gOdFE0J6GSjqsjLor8jM/wqbcENIILCm5DQp3EP8Aod5Jdq
SsVtL1ZkOTHx2lvFu5rCyhoN65bTZ1WkIkpUmOJ7+isPFmFR4DCKvtCHsz6fTJ2VtjfoVi1LlUP8
0fK8Qm6W6F3lKilt9NgHyLL2zXxdqToBLsTQAxRqOODAe1eDB1Px/cXqd0mOksl6tqsxcAgkM/k+
9Nr+O4Gq5LPnqs/C4QGY2dnBfVXZNAECVAlyMQju43e8E7C69jYqISW9sXTyERzN9Gu49Gs3rWUW
oc07taw3+OParb/UkwBsd1Y61wC9yOqg2hqnfZ66+pngbOdDLzOu+GaOnCFkeyKvZGN6bApZQwA2
tr3t4D2tkOeEKLbMKdBrvmwOwEza/X0dxZGXpmrknpAObv+ukB5pLd//f1tqv623CNcA9r93zty/
CO2LmodE1xGtzYNIP2IywaKSvK7Tvv151OMjPw7O41bZdpeDWD2cvc8JvjOvydVga9As5kzHOPgN
MYe2sbEN3rm0JYMhT/CbJ48VuoBBFH7nq1LpSvWCkozzRWXEmcKfm5SLih796jBdxoEr35JJqY5G
+cW9r6S/lqXHd1WArDoA4uortoXEFvFS+UGcd2/dU1eCG3FrZb3PfXdNlY/2fgZ7ii/Q8itnQLq3
6iSqM82lxQXO8Nu0A8D6hUelCTiJ8AjdEbnd/SX1y79/vB1MkSKmGGE3qVKUxRwFsehczUh4rkwe
QgXq48OpA26q1jcZFUgpkb17AIqCt1/0Hx6mduNtdh1zMtqHLGBBdSWwddTdK7VzU6hxsFKouw/b
qpBHdOa5KFZQ4LarPw2xI4TltMAcgUyIhIZfmAnR+nF/A7SnZFspL56oBMcX2yTp6NyLRXvlpnGC
9H5Vg5Bui408cJm+ncCC7pkNtBTaqlrjG7/pIdLAG3s/J8VD5dbQM1TBwF97PlaeXQf/zT8UQUtA
JhDknbwmMSlZbsIpmPeI1PS4Cn27dXVV9bUIU82hRrGbvSf/bNJnXMj07ORW9kKcxoCHRqu+gelH
uE3MLINJ7S/KgGpEf0NbP0SpDuEGM5AYJ/vE4tUygVb0j9T2wEBsoNGYhhSscwr7SqrZeIZgSG6u
/Gt5vhReCaH9fQ5zl0bCg0wu+3RiX4ouIhtoa2q8zBAS5xveSRs9UeMrqFYSsGUhuVujcEv0w81H
cWBjF2z9spQQ2Ia4dIGiOp+1qWov2xrD1QNnNG39lmA/AMvAHpUARInn5dZprfKWBSwJOvk9NPSU
/EHHPSRw6xl6WZWFZXycWLuYMRASflKyxrNNvTBdxt+BGELOYANvSdKC0W4thLvCnIs5XStsLa3P
J4Pyp8vLdGVrEh2Yx5Tuve2Q0HnCEZdfN1c8dnYX0sVbY1WfOxAN+p4q9YBJLr0TN9FgiQTP9QN9
DNLxlucP4CmKMacN1jOROgnfX1Yp6FTWgZ1yCUYRLEGOMbMsoT/vsCEbRLClC7T4+egpoc47Dk2a
o2AkwmpAt424mlRW9yNo9BuEqpcPp4LYBM9KODnmvI8YijhFrjR61QvdQ7vSOjObXSCOaaLKUA5e
h5deUbzSyAhL/4OjfLHDdSVSLpGVg627jIGub7FLxCjPBm0mOrUlSknIZX8051CdrzITuLrzVoen
9SPQr7dPiRGO7NOfGu6I7Pon8uT7GIM8/jDr4L3Jdf9VWOWRXw9+oSvjDdTgMhyTHVqABRjdN727
pEcQ9DtaJKI4AlcbhOSANBBZ0vsxzlpQMvoBBpE46sn6biD/3B80L1Mqfg1/g91knJCXlWQbISuE
cpjH9kNxgL/Sa1bc0gp0KmP+wY3bjdX1A2MZw6nX31cw6FhahDuRkfFswiyu19MpbDZs79DJpG4N
Cqn3VMarC+fFpr02+tgU+iz17twM5HHBuWi48G3RfYPjVKwhFMQ2TBlTp7QBmvHSev+Es3B4nv4T
dBursy3sB6VftFceOvvgYJxSO3uWyEUlgA0c+Zt49LeGqe6scRhSRgh0wLKWsYYDPJJ/Nor/fUzU
Iro3YXBAm2nTqpjwOa6Htb1SNVPOhUfpjfvmGqXYGLnRcX4dcZ4v0eo4DtEUidEOYb/j0ISHt3F1
mM250DByiDxdUui1C2maSCa91JlxedwGAgI1zhCTYCioIfZl9MHhm/dgVDGoESbMSAbLL80PaHvY
7S8/DToefe6Zwuwliy2c+hEIZtrPMWsVQsV9/fgVvuAlz9B7jwemOAm1p2BLcTsWQiUkdOVl46bn
MNLC3pFGV62bjfNb4SIaKLuj0WHnG1ifNEe40p7c6AI3xr1DS+E79rWoeqAigtsWR6uAkrM7A/c/
nxAV+z2qKHLQf3EsRszjiW7NGH9BslX/rOcE/TSFDMtnxkPvuQamZBVJYtUq8bC+aPQuQtXfZVT3
/OcGBuFTJT/d4IXcW6OCfWQ4aywIO98RYwUbgNIyry1qY9G1CzVAe0s7m3Jh88jKAcFX1MJBGbfA
Xa4KGJ8lla8T7XdyP2OObIBKsaL7k9/rQvrVbjob5E3K0mWzFMAR3XYxabF12I4Vj3ZU0YABE/ju
t0Me2Q5My7vWRViMW23kHhnKO0F+e8ZhDidWruz6uBV3+NxKEWFP83SvFUO5AhNqE/qLcHWfQhuk
D8rgch5l7F4l6KiUHOuQkxOAIPDPv9mUkGjaqCL0CgSxwzsOrJKoz1ozmdoZocw0AUltc1wbggve
qSssJ+w4oRl9MKLMcQuAABacSIIyAv0nZq27TlP4FniaSK4dKGOe+DhXU6Zz5S3bEBfEFhj+6D9M
cxKf44FqU7UOxVhNjYh0DzN0t+mNSGlUXHKmORpdLSx7DWcYPeGEeTnW3cQiugeBzthr5L8oSgqj
bvw/5LkfxlSOef0rz8XC759FrzCsHD/BsEpeOgkqLU/pIACXU1zOeGHBqsn5/1g5CmasozyPOSml
7HBQKSEckeWCBljUnT4NiOnEpOqanDbeEi/abQ1MYu3LEsMJYZcc/KdAvc3xNdZ9onlJy1zz+S74
YuDjP0yx3gz01Qe8f219tzG02ldpn/2ua/ynCctRH17lOXxId5KaN2apg1OcUoSGTqLvEMFQMLV2
ZezFYKdcKyoXB9eSTYOA0nE2y+4zU8bNPpQredioiGj0HK2XZHlxiXq7eHeDVCia0N9fy0HeVE1c
HPCwrIdaewWfpvJ0e1IDW4mQ9ZJjSZWwer58bgaePbtQkKEN2GzMeEbz06diSLieGqkIzQ/bBA5S
EGnrqOfrhlKFyf9Ak7lwkB474HlL+I7tsvzKSeQQSxZQ35WFvKl30GEs0jysE0AOzGfo4UPINCsr
9D2bFm2TSxC5Ajw2InRlOM/W8l0W/D2lwHEo0odEACqA17kSS5vIjO0HgNccjEuAwJdOe9uIblMR
idpQ6embrVwgqicguoCZZ2RhYrNhTie9efO06nSoKw9cdo/DUZkcbraDnhEJg9YausF3wuChUCFS
Apleesszi9PDPKLyveMw9OhpMCpSiN5ujHdCTi30zZRCRPszlQgitKIIvoAAc7NTMgzYZUaPRJzQ
d11Uq6Z/w8ziNrtR5g3aJ3WvDIu/ESoVNuGvhBgkyWU2XhCBaiDwkNse8bzbRRsezPgYFmbgOqeo
O0T4f+4WEdxf+dlvy6d8XfWhEHao9NpOvyjuNiVbVgzjSHl63zZ7NjMMdRzOTi3DQuqYNw/59/zT
yoN9VplDlr5VCBxso3nO5NobZeZZi5TaUMQrFFueGj5KammaxluN7DF70icqufnkiURjjfvNlV3d
xWZz1VjiXUgjVMAFGWuYmcZr4CTE0iLWYiN1Zf74PeO1gyCkNcvcmoozZahJogcXomVub7/v3edO
LHgAmAp55kg9ZWHsYVFzVGfltlOkQAXyWu1y93L40gqh5eMJw/iQWB5FM7dhLQPMeSer5V73px3y
iJ4FS/0I6iOVueN/jRPkcaNwlWAMQRJwJASqQODSXfARUKb3Sru9D5aWEGzLQtQgNlKwtbr4KaRl
TqlDzOB/ea7KIk8JCdWK7TNLjtW+ilw0njAWM5/CWdI1XdKifPgwADNVMcP0fDSgnk9+8/uzPpSv
bRObbdYZMvjbzm1RsXGNmIdv/FmCY94LwXiI0yY8Bv7cqfU1S/6lKuev0ke7VIu9TLSaIU8CNY0V
sBDdtbay/1/+ywK/mTaHgcrvSV7s3BBOZWt3jEfi1ELRBZH+FjaBjeIKUiiDuNbama+Pm2MenbaO
2oh+/oCiJqwLXBZ7sW8st34TdT5FNMopCYgEMwEIWMWczwBvv/xp1ekSE+TvTjVzzL9QhDq8TbgS
2YDwDv+YWemmYzhiHDKIIvFu8Z86KMUmx5duCL9PbI61ns0wZLUM1pA4ZxLdC5IsYiqLMXdzti81
FmQ2lq5JU+jVRFYVMQQdQnC8aONkmnjia6MgugNx7/wD19oNd7gfOjfORdHLPp9FqbyLbGT6SrEf
lfK8dg9yDgaXNJQ+RWDD9q3iSAme9LoT1Oc5icZZzW8IWyQnSJyO9jxMKoc7VrDaqeBWBnhQpJ5L
z5GTxv5364qCT7cKXM4eYVzni15l6dKDkNNXEjLUB3E51+vA7VWEh1rLFKHXNqqDMmhzsvRdllJF
my3jcyk4H3jYKQA3RNUQaPniuGipm1xZPKFEqJOnlMWP7lnNZleZvMofzgf/vDDhKbrqvHE3FXqk
gz5TLYdJ0IfKnMVk/xIIMYAP58TU4+S+cT37ettm+zzL9UEHdt8u0zRWGMyJMM0mvJ0b5zSA4dw/
LvtUMlovT3Alnw5ps+OAJI8M3B8haIde+tF9BlmSxh6xojK/hF5CXzyoZSjMu2qz58tWQFOQQEu/
fOJPuwi5OGyI+12ZtO3Gtlifziuj3TEOwOE23juspHQ1iQcn5Hft8uYs7GwGGwxuPmrGc0epXjbQ
cQC2ThkpJVElB7DrOVGvwwBli/8hAulSes6eEOmR47h4SKf/yPTcW539GiWO/O9gHIDiZYiG3Bpq
hSEyVZ4GF1nKvToFIpk6/5Vopykup6K6Ilyas1UtQ4Pp7y8FZjZe049troottssxg7woGd+vB5Eh
IO4t1ht4e/maFZWAyzcAEkDtitSKP2QMdpfPJsejmqsvD5nJAadirrxmhVWE+wZQvuLECZSFkKf7
0Zxe3SFzv6X+MH57XF8ONrCUI8hfhPqM33k8x6pk6K3GJN3wuhdXjpGUzZPi43k83aU5Rag7nSpe
B7XNY97AviFZioDuHf/12hQoqKwy0D6kIgIg5AofdDFDRvHeHB3gcIVCAmJFa8MO4N92Z63YFRMp
w7ICzzLTCqukUGnuJz2jW8rEjrP28aQRWA942rYVIAX9F26gkCWNWhVUNA5y/QQrn8cvoXR3RY2k
JobYnaZVORt3qf9Uc1QzeVFRQlzF3KJgrusEAUezI8WrfM2TLBvGXOjD1G3HSRbbuFt4HPn6g57O
/e5dFm2GZXdiOZ2ebCZ9yyvksQqCkfU1wXrEpecigCJznP2kZO4TH9yp86a/E7tapib8Rw4N5kfc
R8mJGBQMW8beq1j26MexHtH9R8tnoi69iT11P2gVTseD+8/Tv4yJEjOHkwJyKn6APnmdow+UjEE1
qEnCJYyn4xnF+NQyV5jr0R8dvflk8j9Nqh95N8Z6+B/v5EMK2tbbLOBcn7oTUlIrUCC+N0fMl9F3
+YLEuZGydlUJUeo4EzSuIvWG1DL3Z8JhKAaUayeYTItl5XXrm+HSewRzaRHW2lepJ+MQnPx0ty44
aCSt5x1Xx43JWDK5N3lAkupiMe/TuB7SpvoLUREFwriwi9WX6w5kgvicEEbD/mqoWLBaFar15pIu
K7v5CfXkxGXpDhd8j6dauPjK1Z40hKlC9yDKiXvE36l9yYchtBimETVs+fW1A4n6RSoX63o0Njz6
cghxNfDuR8qj+UpnIldgPKk8gVPo1BhIueac84Y7r/pDmkoI80JbzpWPsCXjjrSJF1rXhvox0tgX
pclBYc7+JCrIwBUqOjP7t9yrPj9oSK6zy/w+TAZ3nkZS0LEYJ/6NcmvYA+LJ+fEQqLcDTlPyYijo
bJlNKR3Rn65s7FSKcSa94kJPFsRN8AsdW+7S9imUkJJIuqWl402XTqxG4tURn1QrTIPb2r5q+eX3
eruUEy/K6pQG5+mZ06SNuYVEDxqvwEVaUiHhzuaiXY5k2dtxiIJvaPjZqsN6boflgHXDOa8/nLBz
UiFbQVfXOocbUiTs1C82v0QQjI7m+8NUjRTryub0YUtknY7AMpkYZSyqiYWKGD4OY0tsV5UDvelX
HrzPrAreG2aRrkruimJ/OzXO0k7FpSSgwwLpSvTZ1hYJdcWfMvS7remQ/+OQ6ByQRQX8YYD8J3jM
l/YnaFFaV89sly8AiQ6MPIVc+Y1VPuqA65IiEkMcvxe2HPHSYkhocnpUEeP6dMt2G2VSIpKsqn4B
EPP/nYEO9WV3U+BLZXj3dEwpp/KOaLQB9h+IDkoiFf+4YFa4iRui/6V0z8CCMELMs8zkESa0bCxI
2YTrRPCXKEUrvVQKOdkktQTlAf0950v/zty0Py+TOTHqFuG98VfbtzG84kb1DnyXH3NbpoTCe3FR
+jaGCqWRZB9YbrvOW94G7k6kr/QY6k/W79IrO+FVbBCxd/20WryUbZmfM0dxoIAq9Z2VVCaJbaJf
8L99yN7p2ADCkHb+xsvNQXoIe7d3t13mpd+EzzzHUxQyRWIbUXFKOARGbFjKeilCAGVCsa8O14uw
fjLjqLgQq9nrO92n0rhmz0UIKwleWPsEHmadKKLJzxqZ9D0/Ct8e6EPxgetPOsx60Ni/dsBWQDkY
B5ofivb70AA0qKiB1yNdiv4I7cTs45mrHoJT9nijovrul+6YIGmtApVCHgIY9tjEr9qxHRoLKucQ
FkrCH2Ct71pMUqlxPN9hh8GQxbvvKwcMA/DU2ns1MF2EjaRVelv/PbVfpBSvyAv2bi7EgdgOJCAr
9s3NXA1JAq2ml1cECM8ZXyl94oWWZV5FrVe/qQnJ3es1i/JPCxjcQvxuAOVe/zKOJUGZoPvstJib
CI5wqmuCYzhXYrTGoUy8brNFVO/Ini24CsQ0Bktvl4JrKnSaX+icAR/b+QQ+RaeXRi+4W0WhDZ3x
gkztYT5cYN04hXaPUhZQO3vgkKIi/SRJAXzES9si8hYrQkuJy1FXyYehs5mVX2OO5Bh0NT9/N0N2
u0MUc3YbnUbS56CUM/Lcwg0VgD8bdVJSd7uiZ8aW+KuR+/FlEqRR9q0361Uxp8N0IQcB4oSp+/Qs
15tCYSlAIcdxNJTwexS6eHpCRqi5b/vBstxMGE1FjhlYWKHoH2LkHLz+faAGCYJt+IFeI3NF/EKI
JasuMzn24PD2SfrrKrI5qdOnintdOsVh4nOB8crKGnEDbg/mUmDFeb+E+Wv3sq6Q5LOD56ul+g26
52gHeeJptaPxf9hOmwRAmwd6ngtX/2H84ERZutd5I2+U12OW35/NF9ipEXupbVlknVNpLtscomcs
qZ8oWcIQ7Oc9RTSak3weIUN5OSICbiUrVvtJC7UuZyuSZ4cN0pMVqpgI83a4SxY/Nb8CiF1NDbA3
pF8vwvuvfoPJD34YOivBMdl4/1IjN82HFXqjo6tGX3Hq2gdSJLUMDv2GIIHOQVmTqOLhqBrkI8Ay
GkwAfkJV+iVs44rX31hyWmusixZiQNQgG0qs1/OsNfK0O6R5kzWdDnTNCl8lzkhwTcvGlYtIyb9a
DQcyWnHdpmTSMGts0WkhysaWmwpXCIgqJ0HKLQUjrKf8TTp0S9Xep4sqD97j2VWaYcxhDOVFUoU/
xinfKojy9uvnjvFALg4BXM5O7V4EwxJP00JMX6B7ETThZE0pfmx7VgAWOjUilUndRY+LDXIm4stO
Z6lT9nnLVpNt014XTdwWpPQOiO06is8u11YlkjeirUwZOsepzOGFNpuE14ULkPU225SaD0TrVc2b
yd70uEWn3St8icheO71vFi3Ad/cuJeCUrSiSVStDDwA+AvnSu5kVWGq/N1zkwp/67RwTb8MO7P9f
l7V8GiWUvBNgQF6rhZKZLoLUxxyYi+F/4dW6DkI8aiIiCqf8L2Wroq2ocR26Ndukx/sqckbAVdXL
ksfSe22ey3rP3Qcsg+q5rMAvWUFlR6Wh5Nysymf8bAKS9P1MPfgudnx927Khl4tlRprIE6hUMDkF
wFDv6ITyJpZkYlBXLX9VFjQNY0aJwqAIiPtyhBk56sUmio1R1uK8jiPSITFnOTBuFTG4ORo//dx2
UKuEQHKF3QgdYjDU4/NeR8cnrIjHL1ybYNd1dfdsxzU1XjOD66R7a+Y/w6TKvpVix0G2LsHXS/1+
ZgXItyCCJFPaTIkP8Q0dUFvxisJKSkZcr1fZ3BTNmFoaBHZuIlafy4lpjAkfShK/fSqPO9HjRvJk
TQzED6tNyJ1Jd8llzJ93Z2Lt0dyavjJUiGyJ0ax4AuOUmBR6NvhxDX706RlpscXKWvxD2jWyKIqH
yc5M734BSZfi8KFhA95uTuxVey1jvyHgygo79fLYColm67vSCL3ssfEeHqFdwZOxFtTXiTUmuq+O
d3a9MvbvBFFwbpWMGRq3bIE1DC8Z95JsJWgJVDjdcU1MnXtYMQXQePzUmgGgNkd1f/5so7yKwelU
Xog/EOWeokle6+ThbgvwLYYt0ALIlOTSouOx5u8Hj1CDXYP40gpbgv/0V+s+fYWR3WZwjIwLYsFT
oMWljxfC7YfA4NQiELdMPUtgiZDMNlQNbC+KDku2Ovh4M5eBNv61KUMuhADfUw2PFeFnu5wS0haq
TmpSJlaelDD0G+g8wb9MJVHfIwxI9WRiZSVbrm+4/FMw+P5Is0FvP2wzIm/WAcMNmCe669sPzTkD
eJ0cCeeUpNKwf26W0fXrjMITH9FLjwdmNPqjKrevzsb0g8ivxf/YRdmlY6fvEbyEJkq6lK1XHB5a
R/bzNxjBjpeiTI6YqIgtNWn0e8v06BYPyJynFaqn5btj87z3KJzhCiFpnRsnnRB31C6AeqQ20nMx
VxlZc7ccsqnqKyp5z6ys2AodoeRyu6OdbNFx6hbSmOECIQHLxKS+JgRwUNyB4Zyd+iRMmn1pIyg4
FvtfQGWjnH9oxE7NLj8vM+BZW5ZFSiPkwbMmU/DWwjGA4y18IzsKvyzsKCFkkIP/ZulQwf1cQ9O8
fBRHF8I8vpRoC8G9FK8vHp8QC4O6t8XVPNh5p8BbkBFD6QfDx5RxP5WOSDSmuWljPpm8Xq898OvN
h+Coz4WcZf/b3y82ZjKDBvuZVFIe3LlzQUPJl4o++mVZ0yO6qUr+xe/hku/KTU4ZfVR+M9rf7QJ+
+KQFBG85As0KoY4+sqrSftK2dfDeHXDxHYa/vLr1V5t9J2+8HOgfiZ0PBsO3GlnRXNYBWRIzIOMm
4lrjNSRmuPPpFO4Hs3X8qayiHbsdqKxNt1xgXrq6gOnXBpd51Heo+omalNYAOFEK2LQclg5vYcCH
b5zKyUZos+gp0S8w2tNIQq/2xSGJ6PxSyjKSh7lhkHM58Z0kfIjKsvwBAW+pkcEfM36WaLRNYvCV
3tRiZHkPt8sWEi5QGaC8sT4tZVe/LiNjCkYlaHuWXBtP8haE9aFUOiMdppxbpBSXBAPG1i4LkwQy
pnBJfa6Q5CkIjL1hH+U3WEyngBAzSpKQCwI02tguXMvlFlL+T7rOHEEJCj6COTAQztE1eiaMd8hc
a73sUYKTe2vQJfWCNkc21fA/ofONWXGKT8fJteIJ/GwB
`protect end_protected
