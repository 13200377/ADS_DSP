library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.filter_types.all;

package testBenchFilterIO is

constant numSamples : integer := 1024;
constant test_input_I : int_arr(0 to numSamples-1)(sampleWidth-1 downto 0):= 
(		to_signed(116,sampleWidth),		to_signed(17,sampleWidth),		to_signed(58,sampleWidth),	to_signed(99,sampleWidth),
		to_signed(-1,sampleWidth),		to_signed(99,sampleWidth),		to_signed(58,sampleWidth),	to_signed(16,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(16,sampleWidth),		to_signed(57,sampleWidth),	to_signed(98,sampleWidth),
		to_signed(-1,sampleWidth),		to_signed(98,sampleWidth),		to_signed(57,sampleWidth),	to_signed(16,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(15,sampleWidth),		to_signed(56,sampleWidth),	to_signed(97,sampleWidth),
		to_signed(-2,sampleWidth),		to_signed(97,sampleWidth),		to_signed(55,sampleWidth),	to_signed(14,sampleWidth),
		to_signed(113,sampleWidth),		to_signed(14,sampleWidth),		to_signed(55,sampleWidth),	to_signed(96,sampleWidth),
		to_signed(-4,sampleWidth),		to_signed(95,sampleWidth),		to_signed(54,sampleWidth),	to_signed(12,sampleWidth),
		to_signed(111,sampleWidth),		to_signed(12,sampleWidth),		to_signed(52,sampleWidth),	to_signed(93,sampleWidth),
		to_signed(-6,sampleWidth),		to_signed(93,sampleWidth),		to_signed(51,sampleWidth),	to_signed(10,sampleWidth),
		to_signed(109,sampleWidth),		to_signed(9,sampleWidth),		to_signed(50,sampleWidth),	to_signed(91,sampleWidth),
		to_signed(-9,sampleWidth),		to_signed(90,sampleWidth),		to_signed(48,sampleWidth),	to_signed(7,sampleWidth),
		to_signed(106,sampleWidth),		to_signed(6,sampleWidth),		to_signed(47,sampleWidth),	to_signed(87,sampleWidth),
		to_signed(-12,sampleWidth),		to_signed(86,sampleWidth),		to_signed(45,sampleWidth),	to_signed(3,sampleWidth),
		to_signed(102,sampleWidth),		to_signed(2,sampleWidth),		to_signed(43,sampleWidth),	to_signed(84,sampleWidth),
		to_signed(-16,sampleWidth),		to_signed(83,sampleWidth),		to_signed(41,sampleWidth),	to_signed(-1,sampleWidth),
		to_signed(98,sampleWidth),		to_signed(-2,sampleWidth),		to_signed(39,sampleWidth),	to_signed(79,sampleWidth),
		to_signed(-20,sampleWidth),		to_signed(78,sampleWidth),		to_signed(37,sampleWidth),	to_signed(-5,sampleWidth),
		to_signed(94,sampleWidth),		to_signed(-6,sampleWidth),		to_signed(34,sampleWidth),	to_signed(75,sampleWidth),
		to_signed(-25,sampleWidth),		to_signed(74,sampleWidth),		to_signed(32,sampleWidth),	to_signed(-10,sampleWidth),
		to_signed(89,sampleWidth),		to_signed(-11,sampleWidth),		to_signed(29,sampleWidth),	to_signed(70,sampleWidth),
		to_signed(-30,sampleWidth),		to_signed(69,sampleWidth),		to_signed(27,sampleWidth),	to_signed(-15,sampleWidth),
		to_signed(84,sampleWidth),		to_signed(-16,sampleWidth),		to_signed(24,sampleWidth),	to_signed(65,sampleWidth),
		to_signed(-35,sampleWidth),		to_signed(63,sampleWidth),		to_signed(22,sampleWidth),	to_signed(-20,sampleWidth),
		to_signed(78,sampleWidth),		to_signed(-22,sampleWidth),		to_signed(19,sampleWidth),	to_signed(59,sampleWidth),
		to_signed(-41,sampleWidth),		to_signed(58,sampleWidth),		to_signed(16,sampleWidth),	to_signed(-26,sampleWidth),
		to_signed(73,sampleWidth),		to_signed(-27,sampleWidth),		to_signed(13,sampleWidth),	to_signed(54,sampleWidth),
		to_signed(-46,sampleWidth),		to_signed(52,sampleWidth),		to_signed(10,sampleWidth),	to_signed(-31,sampleWidth),
		to_signed(67,sampleWidth),		to_signed(-33,sampleWidth),		to_signed(8,sampleWidth),	to_signed(48,sampleWidth),
		to_signed(-52,sampleWidth),		to_signed(46,sampleWidth),		to_signed(5,sampleWidth),	to_signed(-37,sampleWidth),
		to_signed(61,sampleWidth),		to_signed(-39,sampleWidth),		to_signed(2,sampleWidth),	to_signed(42,sampleWidth),
		to_signed(-58,sampleWidth),		to_signed(41,sampleWidth),		to_signed(-1,sampleWidth),	to_signed(-43,sampleWidth),
		to_signed(55,sampleWidth),		to_signed(-45,sampleWidth),		to_signed(-4,sampleWidth),	to_signed(36,sampleWidth),
		to_signed(-64,sampleWidth),		to_signed(35,sampleWidth),		to_signed(-7,sampleWidth),	to_signed(-49,sampleWidth),
		to_signed(50,sampleWidth),		to_signed(-50,sampleWidth),		to_signed(-10,sampleWidth),	to_signed(30,sampleWidth),
		to_signed(-70,sampleWidth),		to_signed(29,sampleWidth),		to_signed(-13,sampleWidth),	to_signed(-55,sampleWidth),
		to_signed(44,sampleWidth),		to_signed(-56,sampleWidth),		to_signed(-16,sampleWidth),	to_signed(25,sampleWidth),
		to_signed(-75,sampleWidth),		to_signed(23,sampleWidth),		to_signed(-18,sampleWidth),	to_signed(-60,sampleWidth),
		to_signed(38,sampleWidth),		to_signed(-62,sampleWidth),		to_signed(-21,sampleWidth),	to_signed(19,sampleWidth),
		to_signed(-81,sampleWidth),		to_signed(18,sampleWidth),		to_signed(-24,sampleWidth),	to_signed(-66,sampleWidth),
		to_signed(33,sampleWidth),		to_signed(-67,sampleWidth),		to_signed(-27,sampleWidth),	to_signed(14,sampleWidth),
		to_signed(-86,sampleWidth),		to_signed(13,sampleWidth),		to_signed(-29,sampleWidth),	to_signed(-71,sampleWidth),
		to_signed(28,sampleWidth),		to_signed(-72,sampleWidth),		to_signed(-32,sampleWidth),	to_signed(9,sampleWidth),
		to_signed(-91,sampleWidth),		to_signed(8,sampleWidth),		to_signed(-34,sampleWidth),	to_signed(-76,sampleWidth),
		to_signed(23,sampleWidth),		to_signed(-77,sampleWidth),		to_signed(-36,sampleWidth),	to_signed(4,sampleWidth),
		to_signed(-96,sampleWidth),		to_signed(3,sampleWidth),		to_signed(-39,sampleWidth),	to_signed(-80,sampleWidth),
		to_signed(18,sampleWidth),		to_signed(-81,sampleWidth),		to_signed(-41,sampleWidth),	to_signed(0,sampleWidth),
		to_signed(-100,sampleWidth),		to_signed(-1,sampleWidth),		to_signed(-43,sampleWidth),	to_signed(-85,sampleWidth),
		to_signed(14,sampleWidth),		to_signed(-86,sampleWidth),		to_signed(-45,sampleWidth),	to_signed(-4,sampleWidth),
		to_signed(-104,sampleWidth),		to_signed(-5,sampleWidth),		to_signed(-47,sampleWidth),	to_signed(-88,sampleWidth),
		to_signed(11,sampleWidth),		to_signed(-89,sampleWidth),		to_signed(-48,sampleWidth),	to_signed(-8,sampleWidth),
		to_signed(-107,sampleWidth),		to_signed(-8,sampleWidth),		to_signed(-50,sampleWidth),	to_signed(-92,sampleWidth),
		to_signed(7,sampleWidth),		to_signed(-92,sampleWidth),		to_signed(-51,sampleWidth),	to_signed(-11,sampleWidth),
		to_signed(-110,sampleWidth),		to_signed(-11,sampleWidth),		to_signed(-53,sampleWidth),	to_signed(-94,sampleWidth),
		to_signed(5,sampleWidth),		to_signed(-95,sampleWidth),		to_signed(-54,sampleWidth),	to_signed(-13,sampleWidth),
		to_signed(-113,sampleWidth),		to_signed(-14,sampleWidth),		to_signed(-55,sampleWidth),	to_signed(-97,sampleWidth),
		to_signed(3,sampleWidth),		to_signed(-97,sampleWidth),		to_signed(-56,sampleWidth),	to_signed(-15,sampleWidth),
		to_signed(-115,sampleWidth),		to_signed(-16,sampleWidth),		to_signed(-57,sampleWidth),	to_signed(-98,sampleWidth),
		to_signed(1,sampleWidth),		to_signed(-98,sampleWidth),		to_signed(-58,sampleWidth),	to_signed(-17,sampleWidth),
		to_signed(-116,sampleWidth),		to_signed(-17,sampleWidth),		to_signed(-58,sampleWidth),	to_signed(-99,sampleWidth),
		to_signed(0,sampleWidth),		to_signed(-99,sampleWidth),		to_signed(-58,sampleWidth),	to_signed(-17,sampleWidth),
		to_signed(-117,sampleWidth),		to_signed(-17,sampleWidth),		to_signed(-59,sampleWidth),	to_signed(-100,sampleWidth),
		to_signed(0,sampleWidth),		to_signed(-100,sampleWidth),		to_signed(-59,sampleWidth),	to_signed(-18,sampleWidth),
		to_signed(-117,sampleWidth),		to_signed(-17,sampleWidth),		to_signed(-59,sampleWidth),	to_signed(-100,sampleWidth),
		to_signed(0,sampleWidth),		to_signed(-100,sampleWidth),		to_signed(-58,sampleWidth),	to_signed(-17,sampleWidth),
		to_signed(-116,sampleWidth),		to_signed(-17,sampleWidth),		to_signed(-58,sampleWidth),	to_signed(-99,sampleWidth),
		to_signed(0,sampleWidth),		to_signed(-99,sampleWidth),		to_signed(-58,sampleWidth),	to_signed(-16,sampleWidth),
		to_signed(-115,sampleWidth),		to_signed(-16,sampleWidth),		to_signed(-57,sampleWidth),	to_signed(-98,sampleWidth),
		to_signed(2,sampleWidth),		to_signed(-97,sampleWidth),		to_signed(-56,sampleWidth),	to_signed(-15,sampleWidth),
		to_signed(-114,sampleWidth),		to_signed(-14,sampleWidth),		to_signed(-55,sampleWidth),	to_signed(-96,sampleWidth),
		to_signed(4,sampleWidth),		to_signed(-95,sampleWidth),		to_signed(-54,sampleWidth),	to_signed(-13,sampleWidth),
		to_signed(-112,sampleWidth),		to_signed(-12,sampleWidth),		to_signed(-53,sampleWidth),	to_signed(-94,sampleWidth),
		to_signed(6,sampleWidth),		to_signed(-93,sampleWidth),		to_signed(-51,sampleWidth),	to_signed(-10,sampleWidth),
		to_signed(-109,sampleWidth),		to_signed(-9,sampleWidth),		to_signed(-50,sampleWidth),	to_signed(-91,sampleWidth),
		to_signed(9,sampleWidth),		to_signed(-90,sampleWidth),		to_signed(-48,sampleWidth),	to_signed(-7,sampleWidth),
		to_signed(-106,sampleWidth),		to_signed(-6,sampleWidth),		to_signed(-47,sampleWidth),	to_signed(-87,sampleWidth),
		to_signed(12,sampleWidth),		to_signed(-86,sampleWidth),		to_signed(-45,sampleWidth),	to_signed(-3,sampleWidth),
		to_signed(-102,sampleWidth),		to_signed(-2,sampleWidth),		to_signed(-43,sampleWidth),	to_signed(-84,sampleWidth),
		to_signed(16,sampleWidth),		to_signed(-83,sampleWidth),		to_signed(-41,sampleWidth),	to_signed(1,sampleWidth),
		to_signed(-98,sampleWidth),		to_signed(2,sampleWidth),		to_signed(-39,sampleWidth),	to_signed(-79,sampleWidth),
		to_signed(21,sampleWidth),		to_signed(-78,sampleWidth),		to_signed(-36,sampleWidth),	to_signed(5,sampleWidth),
		to_signed(-93,sampleWidth),		to_signed(6,sampleWidth),		to_signed(-34,sampleWidth),	to_signed(-75,sampleWidth),
		to_signed(25,sampleWidth),		to_signed(-73,sampleWidth),		to_signed(-32,sampleWidth),	to_signed(10,sampleWidth),
		to_signed(-89,sampleWidth),		to_signed(11,sampleWidth),		to_signed(-29,sampleWidth),	to_signed(-70,sampleWidth),
		to_signed(30,sampleWidth),		to_signed(-68,sampleWidth),		to_signed(-27,sampleWidth),	to_signed(15,sampleWidth),
		to_signed(-83,sampleWidth),		to_signed(17,sampleWidth),		to_signed(-24,sampleWidth),	to_signed(-64,sampleWidth),
		to_signed(36,sampleWidth),		to_signed(-63,sampleWidth),		to_signed(-21,sampleWidth),	to_signed(21,sampleWidth),
		to_signed(-78,sampleWidth),		to_signed(22,sampleWidth),		to_signed(-18,sampleWidth),	to_signed(-59,sampleWidth),
		to_signed(41,sampleWidth),		to_signed(-58,sampleWidth),		to_signed(-16,sampleWidth),	to_signed(26,sampleWidth),
		to_signed(-72,sampleWidth),		to_signed(28,sampleWidth),		to_signed(-13,sampleWidth),	to_signed(-53,sampleWidth),
		to_signed(47,sampleWidth),		to_signed(-52,sampleWidth),		to_signed(-10,sampleWidth),	to_signed(32,sampleWidth),
		to_signed(-67,sampleWidth),		to_signed(33,sampleWidth),		to_signed(-7,sampleWidth),	to_signed(-47,sampleWidth),
		to_signed(53,sampleWidth),		to_signed(-46,sampleWidth),		to_signed(-4,sampleWidth),	to_signed(38,sampleWidth),
		to_signed(-61,sampleWidth),		to_signed(39,sampleWidth),		to_signed(-1,sampleWidth),	to_signed(-42,sampleWidth),
		to_signed(58,sampleWidth),		to_signed(-40,sampleWidth),		to_signed(2,sampleWidth),	to_signed(44,sampleWidth),
		to_signed(-55,sampleWidth),		to_signed(45,sampleWidth),		to_signed(5,sampleWidth),	to_signed(-36,sampleWidth),
		to_signed(64,sampleWidth),		to_signed(-34,sampleWidth),		to_signed(8,sampleWidth),	to_signed(49,sampleWidth),
		to_signed(-49,sampleWidth),		to_signed(51,sampleWidth),		to_signed(10,sampleWidth),	to_signed(-30,sampleWidth),
		to_signed(70,sampleWidth),		to_signed(-29,sampleWidth),		to_signed(13,sampleWidth),	to_signed(55,sampleWidth),
		to_signed(-44,sampleWidth),		to_signed(57,sampleWidth),		to_signed(16,sampleWidth),	to_signed(-24,sampleWidth),
		to_signed(76,sampleWidth),		to_signed(-23,sampleWidth),		to_signed(19,sampleWidth),	to_signed(61,sampleWidth),
		to_signed(-38,sampleWidth),		to_signed(62,sampleWidth),		to_signed(22,sampleWidth),	to_signed(-19,sampleWidth),
		to_signed(81,sampleWidth),		to_signed(-18,sampleWidth),		to_signed(24,sampleWidth),	to_signed(66,sampleWidth),
		to_signed(-33,sampleWidth),		to_signed(67,sampleWidth),		to_signed(27,sampleWidth),	to_signed(-14,sampleWidth),
		to_signed(86,sampleWidth),		to_signed(-12,sampleWidth),		to_signed(29,sampleWidth),	to_signed(71,sampleWidth),
		to_signed(-28,sampleWidth),		to_signed(72,sampleWidth),		to_signed(32,sampleWidth),	to_signed(-9,sampleWidth),
		to_signed(91,sampleWidth),		to_signed(-7,sampleWidth),		to_signed(34,sampleWidth),	to_signed(76,sampleWidth),
		to_signed(-23,sampleWidth),		to_signed(77,sampleWidth),		to_signed(37,sampleWidth),	to_signed(-4,sampleWidth),
		to_signed(96,sampleWidth),		to_signed(-3,sampleWidth),		to_signed(39,sampleWidth),	to_signed(80,sampleWidth),
		to_signed(-18,sampleWidth),		to_signed(82,sampleWidth),		to_signed(41,sampleWidth),	to_signed(0,sampleWidth),
		to_signed(100,sampleWidth),		to_signed(1,sampleWidth),		to_signed(43,sampleWidth),	to_signed(85,sampleWidth),
		to_signed(-14,sampleWidth),		to_signed(85,sampleWidth),		to_signed(45,sampleWidth),	to_signed(4,sampleWidth),
		to_signed(104,sampleWidth),		to_signed(5,sampleWidth),		to_signed(47,sampleWidth),	to_signed(88,sampleWidth),
		to_signed(-11,sampleWidth),		to_signed(89,sampleWidth),		to_signed(48,sampleWidth),	to_signed(7,sampleWidth),
		to_signed(107,sampleWidth),		to_signed(8,sampleWidth),		to_signed(50,sampleWidth),	to_signed(91,sampleWidth),
		to_signed(-8,sampleWidth),		to_signed(92,sampleWidth),		to_signed(51,sampleWidth),	to_signed(10,sampleWidth),
		to_signed(110,sampleWidth),		to_signed(11,sampleWidth),		to_signed(52,sampleWidth),	to_signed(94,sampleWidth),
		to_signed(-5,sampleWidth),		to_signed(94,sampleWidth),		to_signed(54,sampleWidth),	to_signed(13,sampleWidth),
		to_signed(112,sampleWidth),		to_signed(13,sampleWidth),		to_signed(55,sampleWidth),	to_signed(96,sampleWidth),
		to_signed(-3,sampleWidth),		to_signed(96,sampleWidth),		to_signed(55,sampleWidth),	to_signed(15,sampleWidth),
		to_signed(114,sampleWidth),		to_signed(15,sampleWidth),		to_signed(56,sampleWidth),	to_signed(97,sampleWidth),
		to_signed(-2,sampleWidth),		to_signed(98,sampleWidth),		to_signed(57,sampleWidth),	to_signed(16,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(16,sampleWidth),		to_signed(57,sampleWidth),	to_signed(98,sampleWidth),
		to_signed(-1,sampleWidth),		to_signed(99,sampleWidth),		to_signed(58,sampleWidth),	to_signed(16,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(16,sampleWidth),		to_signed(58,sampleWidth),	to_signed(99,sampleWidth),
		to_signed(0,sampleWidth),		to_signed(99,sampleWidth),		to_signed(58,sampleWidth),	to_signed(16,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(16,sampleWidth),		to_signed(58,sampleWidth),	to_signed(99,sampleWidth),
		to_signed(-1,sampleWidth),		to_signed(98,sampleWidth),		to_signed(57,sampleWidth),	to_signed(16,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(16,sampleWidth),		to_signed(57,sampleWidth),	to_signed(98,sampleWidth),
		to_signed(-2,sampleWidth),		to_signed(97,sampleWidth),		to_signed(56,sampleWidth),	to_signed(15,sampleWidth),
		to_signed(114,sampleWidth),		to_signed(15,sampleWidth),		to_signed(55,sampleWidth),	to_signed(96,sampleWidth),
		to_signed(-3,sampleWidth),		to_signed(96,sampleWidth),		to_signed(55,sampleWidth),	to_signed(13,sampleWidth),
		to_signed(112,sampleWidth),		to_signed(13,sampleWidth),		to_signed(54,sampleWidth),	to_signed(94,sampleWidth),
		to_signed(-5,sampleWidth),		to_signed(94,sampleWidth),		to_signed(52,sampleWidth),	to_signed(11,sampleWidth),
		to_signed(110,sampleWidth),		to_signed(10,sampleWidth),		to_signed(51,sampleWidth),	to_signed(92,sampleWidth),
		to_signed(-8,sampleWidth),		to_signed(91,sampleWidth),		to_signed(50,sampleWidth),	to_signed(8,sampleWidth),
		to_signed(107,sampleWidth),		to_signed(7,sampleWidth),		to_signed(48,sampleWidth),	to_signed(89,sampleWidth),
		to_signed(-11,sampleWidth),		to_signed(88,sampleWidth),		to_signed(47,sampleWidth),	to_signed(5,sampleWidth),
		to_signed(104,sampleWidth),		to_signed(4,sampleWidth),		to_signed(45,sampleWidth),	to_signed(85,sampleWidth),
		to_signed(-14,sampleWidth),		to_signed(85,sampleWidth),		to_signed(43,sampleWidth),	to_signed(1,sampleWidth),
		to_signed(100,sampleWidth),		to_signed(0,sampleWidth),		to_signed(41,sampleWidth),	to_signed(82,sampleWidth),
		to_signed(-18,sampleWidth),		to_signed(80,sampleWidth),		to_signed(39,sampleWidth),	to_signed(-3,sampleWidth),
		to_signed(96,sampleWidth),		to_signed(-4,sampleWidth),		to_signed(37,sampleWidth),	to_signed(77,sampleWidth),
		to_signed(-23,sampleWidth),		to_signed(76,sampleWidth),		to_signed(34,sampleWidth),	to_signed(-7,sampleWidth),
		to_signed(91,sampleWidth),		to_signed(-9,sampleWidth),		to_signed(32,sampleWidth),	to_signed(72,sampleWidth),
		to_signed(-28,sampleWidth),		to_signed(71,sampleWidth),		to_signed(29,sampleWidth),	to_signed(-12,sampleWidth),
		to_signed(86,sampleWidth),		to_signed(-14,sampleWidth),		to_signed(27,sampleWidth),	to_signed(67,sampleWidth),
		to_signed(-33,sampleWidth),		to_signed(66,sampleWidth),		to_signed(24,sampleWidth),	to_signed(-18,sampleWidth),
		to_signed(81,sampleWidth),		to_signed(-19,sampleWidth),		to_signed(22,sampleWidth),	to_signed(62,sampleWidth),
		to_signed(-38,sampleWidth),		to_signed(61,sampleWidth),		to_signed(19,sampleWidth),	to_signed(-23,sampleWidth),
		to_signed(76,sampleWidth),		to_signed(-24,sampleWidth),		to_signed(16,sampleWidth),	to_signed(57,sampleWidth),
		to_signed(-44,sampleWidth),		to_signed(55,sampleWidth),		to_signed(13,sampleWidth),	to_signed(-29,sampleWidth),
		to_signed(70,sampleWidth),		to_signed(-30,sampleWidth),		to_signed(10,sampleWidth),	to_signed(51,sampleWidth),
		to_signed(-49,sampleWidth),		to_signed(49,sampleWidth),		to_signed(8,sampleWidth),	to_signed(-34,sampleWidth),
		to_signed(64,sampleWidth),		to_signed(-36,sampleWidth),		to_signed(5,sampleWidth),	to_signed(45,sampleWidth),
		to_signed(-55,sampleWidth),		to_signed(44,sampleWidth),		to_signed(2,sampleWidth),	to_signed(-40,sampleWidth),
		to_signed(58,sampleWidth),		to_signed(-42,sampleWidth),		to_signed(-1,sampleWidth),	to_signed(39,sampleWidth),
		to_signed(-61,sampleWidth),		to_signed(38,sampleWidth),		to_signed(-4,sampleWidth),	to_signed(-46,sampleWidth),
		to_signed(53,sampleWidth),		to_signed(-47,sampleWidth),		to_signed(-7,sampleWidth),	to_signed(33,sampleWidth),
		to_signed(-67,sampleWidth),		to_signed(32,sampleWidth),		to_signed(-10,sampleWidth),	to_signed(-52,sampleWidth),
		to_signed(47,sampleWidth),		to_signed(-53,sampleWidth),		to_signed(-13,sampleWidth),	to_signed(28,sampleWidth),
		to_signed(-72,sampleWidth),		to_signed(26,sampleWidth),		to_signed(-16,sampleWidth),	to_signed(-58,sampleWidth),
		to_signed(41,sampleWidth),		to_signed(-59,sampleWidth),		to_signed(-18,sampleWidth),	to_signed(22,sampleWidth),
		to_signed(-78,sampleWidth),		to_signed(21,sampleWidth),		to_signed(-21,sampleWidth),	to_signed(-63,sampleWidth),
		to_signed(36,sampleWidth),		to_signed(-64,sampleWidth),		to_signed(-24,sampleWidth),	to_signed(17,sampleWidth),
		to_signed(-83,sampleWidth),		to_signed(15,sampleWidth),		to_signed(-27,sampleWidth),	to_signed(-68,sampleWidth),
		to_signed(30,sampleWidth),		to_signed(-70,sampleWidth),		to_signed(-29,sampleWidth),	to_signed(11,sampleWidth),
		to_signed(-89,sampleWidth),		to_signed(10,sampleWidth),		to_signed(-32,sampleWidth),	to_signed(-73,sampleWidth),
		to_signed(25,sampleWidth),		to_signed(-75,sampleWidth),		to_signed(-34,sampleWidth),	to_signed(6,sampleWidth),
		to_signed(-93,sampleWidth),		to_signed(5,sampleWidth),		to_signed(-36,sampleWidth),	to_signed(-78,sampleWidth),
		to_signed(21,sampleWidth),		to_signed(-79,sampleWidth),		to_signed(-39,sampleWidth),	to_signed(2,sampleWidth),
		to_signed(-98,sampleWidth),		to_signed(1,sampleWidth),		to_signed(-41,sampleWidth),	to_signed(-83,sampleWidth),
		to_signed(16,sampleWidth),		to_signed(-84,sampleWidth),		to_signed(-43,sampleWidth),	to_signed(-2,sampleWidth),
		to_signed(-102,sampleWidth),		to_signed(-3,sampleWidth),		to_signed(-45,sampleWidth),	to_signed(-86,sampleWidth),
		to_signed(12,sampleWidth),		to_signed(-87,sampleWidth),		to_signed(-47,sampleWidth),	to_signed(-6,sampleWidth),
		to_signed(-106,sampleWidth),		to_signed(-7,sampleWidth),		to_signed(-48,sampleWidth),	to_signed(-90,sampleWidth),
		to_signed(9,sampleWidth),		to_signed(-91,sampleWidth),		to_signed(-50,sampleWidth),	to_signed(-9,sampleWidth),
		to_signed(-109,sampleWidth),		to_signed(-10,sampleWidth),		to_signed(-51,sampleWidth),	to_signed(-93,sampleWidth),
		to_signed(6,sampleWidth),		to_signed(-94,sampleWidth),		to_signed(-53,sampleWidth),	to_signed(-12,sampleWidth),
		to_signed(-112,sampleWidth),		to_signed(-13,sampleWidth),		to_signed(-54,sampleWidth),	to_signed(-95,sampleWidth),
		to_signed(4,sampleWidth),		to_signed(-96,sampleWidth),		to_signed(-55,sampleWidth),	to_signed(-14,sampleWidth),
		to_signed(-114,sampleWidth),		to_signed(-15,sampleWidth),		to_signed(-56,sampleWidth),	to_signed(-97,sampleWidth),
		to_signed(2,sampleWidth),		to_signed(-98,sampleWidth),		to_signed(-57,sampleWidth),	to_signed(-16,sampleWidth),
		to_signed(-115,sampleWidth),		to_signed(-16,sampleWidth),		to_signed(-58,sampleWidth),	to_signed(-99,sampleWidth),
		to_signed(0,sampleWidth),		to_signed(-99,sampleWidth),		to_signed(-58,sampleWidth),	to_signed(-17,sampleWidth),
		to_signed(-116,sampleWidth),		to_signed(-17,sampleWidth),		to_signed(-58,sampleWidth),	to_signed(-100,sampleWidth),
		to_signed(0,sampleWidth),		to_signed(-100,sampleWidth),		to_signed(-59,sampleWidth),	to_signed(-17,sampleWidth),
		to_signed(-117,sampleWidth),		to_signed(-18,sampleWidth),		to_signed(-59,sampleWidth),	to_signed(-100,sampleWidth),
		to_signed(0,sampleWidth),		to_signed(-100,sampleWidth),		to_signed(-59,sampleWidth),	to_signed(-17,sampleWidth),
		to_signed(-117,sampleWidth),		to_signed(-17,sampleWidth),		to_signed(-58,sampleWidth),	to_signed(-99,sampleWidth),
		to_signed(0,sampleWidth),		to_signed(-99,sampleWidth),		to_signed(-58,sampleWidth),	to_signed(-17,sampleWidth),
		to_signed(-116,sampleWidth),		to_signed(-17,sampleWidth),		to_signed(-58,sampleWidth),	to_signed(-98,sampleWidth),
		to_signed(1,sampleWidth),		to_signed(-98,sampleWidth),		to_signed(-57,sampleWidth),	to_signed(-16,sampleWidth),
		to_signed(-115,sampleWidth),		to_signed(-15,sampleWidth),		to_signed(-56,sampleWidth),	to_signed(-97,sampleWidth),
		to_signed(3,sampleWidth),		to_signed(-97,sampleWidth),		to_signed(-55,sampleWidth),	to_signed(-14,sampleWidth),
		to_signed(-113,sampleWidth),		to_signed(-13,sampleWidth),		to_signed(-54,sampleWidth),	to_signed(-95,sampleWidth),
		to_signed(5,sampleWidth),		to_signed(-94,sampleWidth),		to_signed(-53,sampleWidth),	to_signed(-11,sampleWidth),
		to_signed(-110,sampleWidth),		to_signed(-11,sampleWidth),		to_signed(-51,sampleWidth),	to_signed(-92,sampleWidth),
		to_signed(7,sampleWidth),		to_signed(-92,sampleWidth),		to_signed(-50,sampleWidth),	to_signed(-8,sampleWidth),
		to_signed(-107,sampleWidth),		to_signed(-8,sampleWidth),		to_signed(-48,sampleWidth),	to_signed(-89,sampleWidth),
		to_signed(11,sampleWidth),		to_signed(-88,sampleWidth),		to_signed(-47,sampleWidth),	to_signed(-5,sampleWidth),
		to_signed(-104,sampleWidth),		to_signed(-4,sampleWidth),		to_signed(-45,sampleWidth),	to_signed(-86,sampleWidth),
		to_signed(14,sampleWidth),		to_signed(-85,sampleWidth),		to_signed(-43,sampleWidth),	to_signed(-1,sampleWidth),
		to_signed(-100,sampleWidth),		to_signed(0,sampleWidth),		to_signed(-41,sampleWidth),	to_signed(-81,sampleWidth),
		to_signed(18,sampleWidth),		to_signed(-80,sampleWidth),		to_signed(-39,sampleWidth),	to_signed(3,sampleWidth),
		to_signed(-96,sampleWidth),		to_signed(4,sampleWidth),		to_signed(-36,sampleWidth),	to_signed(-77,sampleWidth),
		to_signed(23,sampleWidth),		to_signed(-76,sampleWidth),		to_signed(-34,sampleWidth),	to_signed(8,sampleWidth),
		to_signed(-91,sampleWidth),		to_signed(9,sampleWidth),		to_signed(-32,sampleWidth),	to_signed(-72,sampleWidth),
		to_signed(28,sampleWidth),		to_signed(-71,sampleWidth),		to_signed(-29,sampleWidth),	to_signed(13,sampleWidth),
		to_signed(-86,sampleWidth),		to_signed(14,sampleWidth),		to_signed(-27,sampleWidth),	to_signed(-67,sampleWidth),
		to_signed(33,sampleWidth),		to_signed(-66,sampleWidth),		to_signed(-24,sampleWidth),	to_signed(18,sampleWidth),
		to_signed(-81,sampleWidth),		to_signed(19,sampleWidth),		to_signed(-21,sampleWidth),	to_signed(-62,sampleWidth),
		to_signed(38,sampleWidth),		to_signed(-60,sampleWidth),		to_signed(-18,sampleWidth),	to_signed(23,sampleWidth),
		to_signed(-75,sampleWidth),		to_signed(25,sampleWidth),		to_signed(-16,sampleWidth),	to_signed(-56,sampleWidth),
		to_signed(44,sampleWidth),		to_signed(-55,sampleWidth),		to_signed(-13,sampleWidth),	to_signed(29,sampleWidth),
		to_signed(-70,sampleWidth),		to_signed(30,sampleWidth),		to_signed(-10,sampleWidth),	to_signed(-50,sampleWidth),
		to_signed(50,sampleWidth),		to_signed(-49,sampleWidth),		to_signed(-7,sampleWidth),	to_signed(35,sampleWidth),
		to_signed(-64,sampleWidth),		to_signed(36,sampleWidth),		to_signed(-4,sampleWidth),	to_signed(-45,sampleWidth),
		to_signed(55,sampleWidth),		to_signed(-43,sampleWidth),		to_signed(-1,sampleWidth),	to_signed(41,sampleWidth),
		to_signed(-58,sampleWidth),		to_signed(42,sampleWidth),		to_signed(2,sampleWidth),	to_signed(-39,sampleWidth),
		to_signed(61,sampleWidth),		to_signed(-37,sampleWidth),		to_signed(5,sampleWidth),	to_signed(46,sampleWidth),
		to_signed(-52,sampleWidth),		to_signed(48,sampleWidth),		to_signed(8,sampleWidth),	to_signed(-33,sampleWidth),
		to_signed(67,sampleWidth),		to_signed(-31,sampleWidth),		to_signed(10,sampleWidth),	to_signed(52,sampleWidth),
		to_signed(-46,sampleWidth),		to_signed(54,sampleWidth),		to_signed(13,sampleWidth),	to_signed(-27,sampleWidth),
		to_signed(73,sampleWidth),		to_signed(-26,sampleWidth),		to_signed(16,sampleWidth),	to_signed(58,sampleWidth),
		to_signed(-41,sampleWidth),		to_signed(59,sampleWidth),		to_signed(19,sampleWidth),	to_signed(-22,sampleWidth),
		to_signed(78,sampleWidth),		to_signed(-20,sampleWidth),		to_signed(22,sampleWidth),	to_signed(63,sampleWidth),
		to_signed(-35,sampleWidth),		to_signed(65,sampleWidth),		to_signed(24,sampleWidth),	to_signed(-16,sampleWidth),
		to_signed(84,sampleWidth),		to_signed(-15,sampleWidth),		to_signed(27,sampleWidth),	to_signed(69,sampleWidth),
		to_signed(-30,sampleWidth),		to_signed(70,sampleWidth),		to_signed(29,sampleWidth),	to_signed(-11,sampleWidth),
		to_signed(89,sampleWidth),		to_signed(-10,sampleWidth),		to_signed(32,sampleWidth),	to_signed(74,sampleWidth),
		to_signed(-25,sampleWidth),		to_signed(75,sampleWidth),		to_signed(34,sampleWidth),	to_signed(-6,sampleWidth),
		to_signed(94,sampleWidth),		to_signed(-5,sampleWidth),		to_signed(37,sampleWidth),	to_signed(78,sampleWidth),
		to_signed(-20,sampleWidth),		to_signed(79,sampleWidth),		to_signed(39,sampleWidth),	to_signed(-2,sampleWidth),
		to_signed(98,sampleWidth),		to_signed(-1,sampleWidth),		to_signed(41,sampleWidth),	to_signed(83,sampleWidth),
		to_signed(-16,sampleWidth),		to_signed(84,sampleWidth),		to_signed(43,sampleWidth),	to_signed(2,sampleWidth),
		to_signed(102,sampleWidth),		to_signed(3,sampleWidth),		to_signed(45,sampleWidth),	to_signed(86,sampleWidth),
		to_signed(-12,sampleWidth),		to_signed(87,sampleWidth),		to_signed(47,sampleWidth),	to_signed(6,sampleWidth),
		to_signed(106,sampleWidth),		to_signed(7,sampleWidth),		to_signed(48,sampleWidth),	to_signed(90,sampleWidth),
		to_signed(-9,sampleWidth),		to_signed(91,sampleWidth),		to_signed(50,sampleWidth),	to_signed(9,sampleWidth),
		to_signed(109,sampleWidth),		to_signed(10,sampleWidth),		to_signed(51,sampleWidth),	to_signed(93,sampleWidth),
		to_signed(-6,sampleWidth),		to_signed(93,sampleWidth),		to_signed(52,sampleWidth),	to_signed(12,sampleWidth),
		to_signed(111,sampleWidth),		to_signed(12,sampleWidth),		to_signed(54,sampleWidth),	to_signed(95,sampleWidth),
		to_signed(-4,sampleWidth),		to_signed(96,sampleWidth),		to_signed(55,sampleWidth),	to_signed(14,sampleWidth),
		to_signed(113,sampleWidth),		to_signed(14,sampleWidth),		to_signed(55,sampleWidth),	to_signed(97,sampleWidth),
		to_signed(-2,sampleWidth),		to_signed(97,sampleWidth),		to_signed(56,sampleWidth),	to_signed(15,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(16,sampleWidth),		to_signed(57,sampleWidth),	to_signed(98,sampleWidth),
		to_signed(-1,sampleWidth),		to_signed(98,sampleWidth),		to_signed(57,sampleWidth),	to_signed(16,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(16,sampleWidth),		to_signed(58,sampleWidth),	to_signed(99,sampleWidth),
		to_signed(-1,sampleWidth),		to_signed(99,sampleWidth),		to_signed(58,sampleWidth),	to_signed(17,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(17,sampleWidth),		to_signed(58,sampleWidth),	to_signed(99,sampleWidth),
		to_signed(-1,sampleWidth),		to_signed(99,sampleWidth),		to_signed(58,sampleWidth),	to_signed(16,sampleWidth),
		to_signed(116,sampleWidth),		to_signed(16,sampleWidth),		to_signed(57,sampleWidth),	to_signed(98,sampleWidth),
		to_signed(-1,sampleWidth),		to_signed(98,sampleWidth),		to_signed(57,sampleWidth),	to_signed(16,sampleWidth),
		to_signed(115,sampleWidth),		to_signed(15,sampleWidth),		to_signed(56,sampleWidth),	to_signed(97,sampleWidth),
		to_signed(-2,sampleWidth),		to_signed(97,sampleWidth),		to_signed(55,sampleWidth),	to_signed(14,sampleWidth) );

constant test_output_I : int_arr(0 to numSamples/phaseCount -1)(sampleWidth-1 downto 0):= 
(		to_signed(19,sampleWidth),		to_signed(55,sampleWidth),		to_signed(98,sampleWidth),	to_signed(87,sampleWidth),
		to_signed(97,sampleWidth),		to_signed(85,sampleWidth),		to_signed(95,sampleWidth),	to_signed(83,sampleWidth),
		to_signed(93,sampleWidth),		to_signed(80,sampleWidth),		to_signed(89,sampleWidth),	to_signed(76,sampleWidth),
		to_signed(85,sampleWidth),		to_signed(71,sampleWidth),		to_signed(79,sampleWidth),	to_signed(65,sampleWidth),
		to_signed(73,sampleWidth),		to_signed(58,sampleWidth),		to_signed(66,sampleWidth),	to_signed(51,sampleWidth),
		to_signed(59,sampleWidth),		to_signed(43,sampleWidth),		to_signed(50,sampleWidth),	to_signed(35,sampleWidth),
		to_signed(42,sampleWidth),		to_signed(26,sampleWidth),		to_signed(33,sampleWidth),	to_signed(17,sampleWidth),
		to_signed(24,sampleWidth),		to_signed(8,sampleWidth),		to_signed(15,sampleWidth),	to_signed(-1,sampleWidth),
		to_signed(5,sampleWidth),		to_signed(-11,sampleWidth),		to_signed(-4,sampleWidth),	to_signed(-20,sampleWidth),
		to_signed(-14,sampleWidth),		to_signed(-29,sampleWidth),		to_signed(-23,sampleWidth),	to_signed(-38,sampleWidth),
		to_signed(-32,sampleWidth),		to_signed(-47,sampleWidth),		to_signed(-40,sampleWidth),	to_signed(-55,sampleWidth),
		to_signed(-48,sampleWidth),		to_signed(-63,sampleWidth),		to_signed(-56,sampleWidth),	to_signed(-71,sampleWidth),
		to_signed(-63,sampleWidth),		to_signed(-77,sampleWidth),		to_signed(-69,sampleWidth),	to_signed(-83,sampleWidth),
		to_signed(-74,sampleWidth),		to_signed(-88,sampleWidth),		to_signed(-79,sampleWidth),	to_signed(-92,sampleWidth),
		to_signed(-83,sampleWidth),		to_signed(-96,sampleWidth),		to_signed(-86,sampleWidth),	to_signed(-99,sampleWidth),
		to_signed(-88,sampleWidth),		to_signed(-100,sampleWidth),		to_signed(-89,sampleWidth),	to_signed(-101,sampleWidth),
		to_signed(-90,sampleWidth),		to_signed(-101,sampleWidth),		to_signed(-89,sampleWidth),	to_signed(-99,sampleWidth),
		to_signed(-87,sampleWidth),		to_signed(-97,sampleWidth),		to_signed(-85,sampleWidth),	to_signed(-94,sampleWidth),
		to_signed(-81,sampleWidth),		to_signed(-90,sampleWidth),		to_signed(-77,sampleWidth),	to_signed(-86,sampleWidth),
		to_signed(-72,sampleWidth),		to_signed(-80,sampleWidth),		to_signed(-66,sampleWidth),	to_signed(-74,sampleWidth),
		to_signed(-59,sampleWidth),		to_signed(-66,sampleWidth),		to_signed(-52,sampleWidth),	to_signed(-59,sampleWidth),
		to_signed(-44,sampleWidth),		to_signed(-51,sampleWidth),		to_signed(-35,sampleWidth),	to_signed(-42,sampleWidth),
		to_signed(-27,sampleWidth),		to_signed(-33,sampleWidth),		to_signed(-18,sampleWidth),	to_signed(-24,sampleWidth),
		to_signed(-8,sampleWidth),		to_signed(-15,sampleWidth),		to_signed(1,sampleWidth),	to_signed(-5,sampleWidth),
		to_signed(11,sampleWidth),		to_signed(4,sampleWidth),		to_signed(20,sampleWidth),	to_signed(13,sampleWidth),
		to_signed(29,sampleWidth),		to_signed(23,sampleWidth),		to_signed(38,sampleWidth),	to_signed(31,sampleWidth),
		to_signed(46,sampleWidth),		to_signed(39,sampleWidth),		to_signed(55,sampleWidth),	to_signed(47,sampleWidth),
		to_signed(63,sampleWidth),		to_signed(55,sampleWidth),		to_signed(70,sampleWidth),	to_signed(62,sampleWidth),
		to_signed(76,sampleWidth),		to_signed(68,sampleWidth),		to_signed(82,sampleWidth),	to_signed(73,sampleWidth),
		to_signed(87,sampleWidth),		to_signed(78,sampleWidth),		to_signed(91,sampleWidth),	to_signed(81,sampleWidth),
		to_signed(94,sampleWidth),		to_signed(84,sampleWidth),		to_signed(96,sampleWidth),	to_signed(86,sampleWidth),
		to_signed(98,sampleWidth),		to_signed(87,sampleWidth),		to_signed(98,sampleWidth),	to_signed(87,sampleWidth),
		to_signed(98,sampleWidth),		to_signed(86,sampleWidth),		to_signed(96,sampleWidth),	to_signed(84,sampleWidth),
		to_signed(94,sampleWidth),		to_signed(81,sampleWidth),		to_signed(91,sampleWidth),	to_signed(77,sampleWidth),
		to_signed(86,sampleWidth),		to_signed(73,sampleWidth),		to_signed(81,sampleWidth),	to_signed(68,sampleWidth),
		to_signed(76,sampleWidth),		to_signed(62,sampleWidth),		to_signed(69,sampleWidth),	to_signed(55,sampleWidth),
		to_signed(62,sampleWidth),		to_signed(47,sampleWidth),		to_signed(54,sampleWidth),	to_signed(39,sampleWidth),
		to_signed(46,sampleWidth),		to_signed(31,sampleWidth),		to_signed(38,sampleWidth),	to_signed(22,sampleWidth),
		to_signed(29,sampleWidth),		to_signed(13,sampleWidth),		to_signed(19,sampleWidth),	to_signed(4,sampleWidth),
		to_signed(10,sampleWidth),		to_signed(-6,sampleWidth),		to_signed(0,sampleWidth),	to_signed(-15,sampleWidth),
		to_signed(-9,sampleWidth),		to_signed(-25,sampleWidth),		to_signed(-18,sampleWidth),	to_signed(-34,sampleWidth),
		to_signed(-27,sampleWidth),		to_signed(-42,sampleWidth),		to_signed(-36,sampleWidth),	to_signed(-51,sampleWidth),
		to_signed(-45,sampleWidth),		to_signed(-60,sampleWidth),		to_signed(-52,sampleWidth),	to_signed(-67,sampleWidth),
		to_signed(-59,sampleWidth),		to_signed(-74,sampleWidth),		to_signed(-66,sampleWidth),	to_signed(-80,sampleWidth),
		to_signed(-72,sampleWidth),		to_signed(-86,sampleWidth),		to_signed(-77,sampleWidth),	to_signed(-91,sampleWidth),
		to_signed(-81,sampleWidth),		to_signed(-94,sampleWidth),		to_signed(-85,sampleWidth),	to_signed(-97,sampleWidth),
		to_signed(-87,sampleWidth),		to_signed(-100,sampleWidth),		to_signed(-89,sampleWidth),	to_signed(-101,sampleWidth),
		to_signed(-90,sampleWidth),		to_signed(-101,sampleWidth),		to_signed(-89,sampleWidth),	to_signed(-100,sampleWidth),
		to_signed(-88,sampleWidth),		to_signed(-99,sampleWidth),		to_signed(-86,sampleWidth),	to_signed(-96,sampleWidth),
		to_signed(-83,sampleWidth),		to_signed(-92,sampleWidth),		to_signed(-79,sampleWidth),	to_signed(-88,sampleWidth),
		to_signed(-74,sampleWidth),		to_signed(-83,sampleWidth),		to_signed(-69,sampleWidth),	to_signed(-77,sampleWidth),
		to_signed(-62,sampleWidth),		to_signed(-70,sampleWidth),		to_signed(-56,sampleWidth),	to_signed(-63,sampleWidth),
		to_signed(-48,sampleWidth),		to_signed(-55,sampleWidth),		to_signed(-40,sampleWidth),	to_signed(-47,sampleWidth),
		to_signed(-31,sampleWidth),		to_signed(-38,sampleWidth),		to_signed(-22,sampleWidth),	to_signed(-29,sampleWidth),
		to_signed(-13,sampleWidth),		to_signed(-20,sampleWidth),		to_signed(-4,sampleWidth),	to_signed(-10,sampleWidth),
		to_signed(6,sampleWidth),		to_signed(-1,sampleWidth),		to_signed(15,sampleWidth),	to_signed(9,sampleWidth),
		to_signed(24,sampleWidth),		to_signed(18,sampleWidth),		to_signed(33,sampleWidth),	to_signed(27,sampleWidth),
		to_signed(42,sampleWidth),		to_signed(36,sampleWidth),		to_signed(51,sampleWidth),	to_signed(44,sampleWidth),
		to_signed(59,sampleWidth),		to_signed(52,sampleWidth),		to_signed(66,sampleWidth),	to_signed(59,sampleWidth),
		to_signed(73,sampleWidth),		to_signed(65,sampleWidth),		to_signed(79,sampleWidth),	to_signed(71,sampleWidth),
		to_signed(85,sampleWidth),		to_signed(76,sampleWidth),		to_signed(89,sampleWidth),	to_signed(80,sampleWidth),
		to_signed(93,sampleWidth),		to_signed(83,sampleWidth),		to_signed(95,sampleWidth),	to_signed(85,sampleWidth),
		to_signed(97,sampleWidth),		to_signed(87,sampleWidth),		to_signed(99,sampleWidth),	to_signed(87,sampleWidth),
		to_signed(98,sampleWidth),		to_signed(87,sampleWidth),		to_signed(97,sampleWidth),	to_signed(85,sampleWidth) );

end package;