-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
XIm1Cv3ZoU+ox/2U5WcLHsLO+V4k8tSR1R1buMECfmtxJ0WfkIbUc8KumHOJA539AvKdwA16ppiU
lbPv8yhp0zGUhj92C1n04EDOBwiEdKhAyh7OYw27C/NBJ7COvcnll/lznNTSISH9gl3DtSv0EuIS
dzQX43Gd5RwabARTny+mZ0sCx/vmXhzlTLvCtV/oGj1Qi/Te4msy50HvfWtVWuv3eETDEeQkGLhy
8DN308WwYU5n+YZRKtxsgdXZrkQS8X2RD5cIkTOB73xoJZGHGVIMZk9ffZL7umdMGeRWv2qQd5X/
/zkx1XWsmRbmoabPDOaO5ApIQM78TrHiufjmNA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 18800)
`protect data_block
ncT8iSn0R2865lZ4vFtLSI5a8hoFEc1bgW3qRCV3pL4gyN8QdIRuo/kDJZqj9UiN/ugjC3wBze0+
R+0vebhnH5qPawRjOiv8/bcMR9KLqumBYgu4BWaLlqy+fjGMBFbXlRO2/XvNbaLcIdMp682arYoU
pfxj2HwFlZgRcHfuuejnhHuOZM8I06N0Zyt5O+x/jybDItAilKGXulh4MkLTbXFGqOrg2GeylfaQ
m6yA8dKYEbMpjscNOC7D4266onil4NAEaEDV94iL4/1u4W+VasfnbNC67Q9xE9fjVtHTxRpwSFk/
86x+WZeFoqPOgdvgpyTg4ydH//HxpTZS+x75CNw5o/1hlxk1E20vvRsxXTQTC57tET58qOj85FUY
tyrFVPFlgq5P0689Uqhw5KkHcNTF5vPte38joA6ThMIWmmcynHjD8rT5t3vq+lR22QdC9eFpsDsb
d1PQGeF3gqa/Ud661EcRPP/5ZmDYmTZySPn8veRz7JXN59g6HjNyKoM2TKeJDc+JspDUAj1UvYVp
cDrCi5f9KjrMK9A22VSgYfRHCr321vXdjr8PO79o08d+OWCYVMm0+RPazTVFeaCMj+H2LD1Heilc
224VAKhBMeumopk4hAHdfmTMdyglB0KVEgukLIzXbk+XjYYsbGBbYM+jE6SOKNk3qKelIIkzjAwd
Zx5aZQQ/Qf/73UXoXK0e9veFEP4Mf5kwCGDPtxqK0OP/06e/jpegwHtkn2nd3GlStO22kmtfL7sW
jqpivCoSdDjeOzKHcuf0Qp+Wwt02IQO1rTDJeoVo0GP+g/mBIgFhrJrCATF2sWlrY71RHhkHnaeU
vOSzzvdxSEC/ucIXiBnMdAfneKwUy0WLCP6rcaXBVb+LppjnAiCKhrw4shir4GajREaGQHmlAh6z
AMMeuQTVSbRd6WT16o81vqPyFPNwPIWWoPC7as0asNnyVAKJWc5L1Rm9w78BYvn3oJ/9llPQkqCo
euvRwqAMeAIoh3rSYuL/J6Krfg5+5pLQycz0MibGSo1PwBZ7cCnfccwUVxA3wFUBetoq3q52uon/
10iRE9CdfU5MzrqETXpvV+QwlVrbFwNn9OQ62TOnQZQsMFZ2ovyd0jyful/T1GogWqhNcSHLtXcm
KPeyX0k1qnulSYI8uvu827tWgyoaskZx5Ww2SsEZRkEOJcy3uYyCTB4/hT2I7yTLWyP67XednYEI
RrbzXTc0Hp3bbZ45hCR/G0Y1mRAJtwkcQFNi6sHwRYQlnaz5de2uuSnNfQ3IXTDeEv0gzrLc1L9+
/jYixiI4LiU7+n9U2cmKYMQBu/EJlKdMqXjlQ8Iqie56MyYlKCSXWytnsGkIuOb5RPw7Nq/wo9w9
8A3rlumKCN9gBiXGs2MBILeaO8iJIfsBgi2hvhgP+CAHb0P9N/thFaszmRoLaDPqB8MLULl3DzBa
crYenkhAWM+JN95YMlZea9/0TqNSiFbv3fGdieeAyMCZfJaYB+Hi8o3SBO+cjreo+0SQTLsXCJlf
0inxwBclVgF4V5NjBKzGTXqK7eTupHB2F91rwlt55Xb2bWSRVspU3i0IFR8+sq6EDPIpSVF32AOr
NNG/nruEQbwdFvh9XZjrXuTOfgqnJG+6YMtbw2bNHKs6Mi8t1b1hQ0TRLfPgUy3ZCSfqGuIUb7Sx
19v25zWKiB9CxExfHrDIibW1+jseZjzPhzjWr6D1IJYzalSMhptsR3CO4Hjd5UfpLvIp09bK2Tvl
PzAZjVwCsUAiLqROgu4AzeT9Fp4BgFWhnVIFvPEq3p/uhYfPDgOJLHEilhGpcbdpsNReNhxyF6Qo
NhnuWvzz19f+bTMBr3dQN5CF7WK75tFFKpH15OFtdKX6hlDacUvYflKsOMPvqqjQ5btxZeNhgudq
sKHA8h+dGG1AVLFCCRKrMcbFjlhYZRRGGVvUS/D7sl2pRZejW2LmqMdemLOFarHoT6pedQCiDqHC
8oIwtn71PQ3DulzsJ3oOuWsn09fb91ogkYUIUmZLqrL8kSXxtycxDTiXr92ljshp23vduwTwi2Nu
l0fFH6qSRSf0Z6hO2ggjO2GCvmzBhYNGlU56Ttw40blRZWMri7HyvjTfxHCXIjR1sZ/Qor6nzqsb
KCLWcFk3/sQBtJL9gJQCyaALNoENiuPHumf4/VGQ4qTuGFfcMilsuVYIIbbasRmjCYe1mDxbQ8s5
VCKFllizFrxlt0NDudyLnSRvAXRb5FYJoQtus3Ed2S3jpsRLPILWdDoQsJChT14mPeWRsuQ9HlbJ
xik1KzGNsX4UXKHSYi7I5Agx+kaPZf+LpsmiM9B26tlowTirUjJIWJ4I0qqII6Hvxgum6MDvUiLZ
xh82XJ1KR4aFKTP33+AzktSn2DGoEhXIVTwV2VTZFuLn9IZIzkLRpiQ63IQzQnOZVX3/Lix/PH0k
kJBZOV+blvGsL/Fg6nmwNLD0H8UJ51aUfhzaiDD0fBLlnF+kMRJqQ33qGuyZAJVx3JOEBm+6dA5j
GufTlB2QuTQ42aVZ0r8pO0wJGv/UPAmLrNTuFN3ffoJ86vUIWhBUCfVfjCAizQawhaVveKGTO4Vm
N0sluin9M9e3kQJfcVvidS8wN0LfIeL/0pNQO7wkv15kmzpb71bEiX7e4tFglp9UG9K5AedtNWot
V4k/qL9d1B4Q484fYNF9nFq+Ncnj6o/ap9F7oCIOlVq4oHQhHiUtBKs81qekpDTz0TsjovK5ctkK
yD+LhovmQ/oG8LPHK+f5AXIuZoFduJOn8qcTOJx47XxEr1Oed9PnENpFHrmg4EyLhV558++W/+Z7
jNvYOP3Vw68xyJg9C4SuZSCJw+RMZkDPL5Nl0tSOGsQip54SBK9V7D+vzPKiqy5Mj1u4zWfFzLq/
F10kTN1iC8dYOUnpB9GHAJLYCza+lDakQtaIW9F1xxh6MsUj94zm2WGhoBjVa8MsIS0rQNNHCJyO
1agncLgewHFI84oXHW09VF+ZZxvqE1olL9fYD5gmWHNovBscI3OxURS+8qK+1fK0RQBtj9QadR6R
JTGHw3czrlruOosYrjFBYbxWMe7bTcvzIHMAEM+fk4BWTWCFUXEOLiE2h/C3EIbC7pdAdLQ9hPXD
ta3PDqcw0ZC8sXWoXmG1V5AjHpjvx6LqLATPtrm1NJBiTLTaYfKPp/56H+xtz/nV3VJif44oUdE7
FmK+X1tE3b8kPZgrm8dlhYuGEthi4kg0BNB90+hHtE5zPlfbZACjygs2rn0PuTFbdtwsv8pTkjJk
FU7/MG/MBqmVIV2uVIxfg3S3/KGTYKrjBHKXS4ZT/kfL1UrWvy8EHEseENUI1yDnwhigi9Pkva6h
zJ/fXCmSHc7RDFgJbzEcPPYdMVFfT8Lna+sw12PXF3n9yc7lsoH6DeWp8Pg0LFJ4gTg01Wd+bv8p
ITYQ97w6jswxinePOV95qqcr2qPLnkOExKC+L2UWWm+GEpJAOyyPuT/PHiiPPruvmCmf17CAZflr
BOMRCOVTLVavNW9wJujGHMNbvYgULoGZOj1p//p2KWQ0lLvAuR6CSmeADIPJN872qY/Z5clqVUsJ
5am/Ctac7G1bDBHfGbukK8IsSv5lMYplKT3mqmFi3qIIZTjUqfeFCxfHedk+2oybMj9nY0Qcm9D1
tJJr11qa1f1rfQkjyENIDTxCT1AHr9bB51bnj7RqNoUVr9DX0MjaxuE6uILb/t4hJjYLsgfMsgae
ZWsDq1sCOIsKfi7S3qatIDfSasr3EWxCIjYFHoE3cEgV7kW4S3OvG6GTXE7Yj2k2yMWuA9dLGKbs
Qy9hqxg21UGR/Tf3RX6WhXjdWKtYmrfAYyez4kPmDM6+kwUutICr408/rXpM8XcVwnWgmTO+UVQF
Q9c/mbU25Bn/gm4UxOb1DHWouUcCERAZIt/cYQBwS/ucYTx911PDPH6grKu/AuiQckFFaxpAwacq
SqjUn4zGvcjT886p80eAnu4Qlk2zdjZ0ocqSa9Qp58GxE6Dn3whzxIEoG4izwzrxvaetaGGm/5A3
/vQ4o1UOPHLPH6vcs7zgRAw6e2/5cC/xBk1bAAREr4tupkL2kXOmwfpxqvVpnABkkVpTpDqG3bCM
/nhkges1LML0c3mwAwicEzUOcWY/yWtDetmlThHTXqfZNjUuyLK9KZT0iXWWOl59npiO5Vn96qCN
ALYK6ReRGE/j0iGm9RKalKovNQh/yXVaW28vI5fzO/mMcTOw/l2tubBLGSeWx9fzcPqbBwrCbUL0
FpBx4ZESEmMvb4pFSEeJ+8DVzyEKIHnJ7JoytcHSn/ytZ7XJOxeEP/lcH8dhidUpOliDcTn8s8uV
JMelko0EiA6vTz2t249L8URbadfQu1i66ARlHxUi4grAhqiwKKmlQRkun/QoLASTzWeSg4plIRYR
6pO4re9b7itpxrkHMs0cx4cbJxqwiOs8s8Xc/tOOvU2Egg4Ob4ElhCnGJcGMIaPpxi8nFu+/IVzf
7r2pDIRVn9qcVN2k2sBpQ3aibRXQm3N3sBLIt3Hwr0e4i1nLrU/Fz9HvL2gFcmLWIsDl1ceBMVKM
eAyV+WiH2UB2Y+c/pQ9eW/GIC5pzC7Pv5WGw9RJwvGNSG6W7/1m8d689oz4plwBzgwjtxJuRmVIU
4s4Se1CIjirduWf2HEXxpgWch5IYUvbzFBuJqjVixIl5JU5sTcM2c61cFwNT7Rm3bR50Cmtjmt6b
OATO+n+ChLHHTsRYQbNtfE1ZVekvw5rscPDo1UP93rudHA2AW0Vf7GbPUoxrs6FiljHaP8GkTeut
yvOPTaVUgc0buuQKAzpif5Bsp8T7gckkTd75V5nUlr28raDTxIFtnETtPrWYBDI2PWnHLsF17PjD
8tlpXbDnDWF0PSququg73bgfKU7zSQYR0bA8KSwMSzNdEUm4mTjKTE3iwIf8znZECtHDJUtzZdB3
SwBGUbn6j6rTWuoE6njoVeHs4TUyoWxUB5RsH63Zg+LT1poluNrYy+W5FPgrbqSuWeTWLtjc2rEb
osKLepsqj0UA4++KBL2Z6uUw7+D+d8DNVcz8d87kx7zjHeQi29sSZZQzcOFZWR+K/QCJrlScFpn6
FSy5hmjrFVb3vj7oOtIxDmW2sMRKDs47+mbBAwFCilQlwIzqoQ1OSl9t8gG+Mk3DH81qyVyvNeTC
k8PUuabshPew6b+nnUq5mhS/3il6SvNSrFHFzoRWu1HBYCdMqzGLKMCRGO/MBXkReh3EeomEdkWz
ba08FOT6+AYBVivjlgC+vT4ASDQM35tQ1hvjMF7R61zcsUWWp8/sp/vzalkUTgrV63ZuWw1fNbDe
9PY/uiONPOucG4EHGhBg++YJLgr8v3g8aZXOeWEV4BLtZstgbRwSQbOsho7A6f3thcJ6U0KszR5E
bdrYtP5S1whSI2e55l00Q/JQOJtVRhLmeUiwpb7kXhm20HNdxffR8pW8B3OVYderHphR62ib2WX4
d9gpLzTLsK4Iu7XlRUPkXSfQP/oT0ON26V9WrSBNY2t5wzj9xB3zhOf1KLaSYWYiC/lucxkcj4O9
YxttPZLDBNyKJJzKHmGlmVU+bPf33GDsGmM6FoyNgiy6M2vdkdU6NIVPh8EfGumyZymBVVokrp4q
5aQJ4B+BrFA9C6cdncPHFrEK4uAJmohS54nqur3x5nU2QNrEV91TxAfDrq2Mi7mvGBurXwycsh0L
ENt5obDDCNkEqlu7uypUWNN8c81CFZmtxA9k4ASBsU/WCI1e0laJTCE0New/u8hHU8HLBwb3t3QC
Grtx6v4LTUClcGtDPsemVh4uLMpzpqjRoKUWC+ttaEgLlxJ8RuGEezfvjfyxhQ3cH2IfRMNpnQCF
XUJkVNjSu1EZ8yp2+sjyq7UZh35GhTW9UDXxBmtM2uLtkxNGAZ1Z2ibKwCavuB2lxdwowi7Smcl2
+wcqFT0JGr67K/pAJVHVDL+HbOz/dOHRtdVZaHWk+139Njt6XTLgZOd/z/gENufsoIyaC9PTCtRX
dQ/OitzoFPPm6YwrhXNwDA+wmfX88BC1Sxhnq1/Eu2pBotcDUl3DUdShDYgCKmSYuzsPN/WPa3iH
ej4wjRjn9++ywSsfoR5ww5Gzsb3y0z7OGs7W7I8cp/ugTgCp5rs1RLoldZSOlBDGDmnzvHaHJ1FP
/m5EKkMBTwlDPV1X4UjxqsR/aZjoSrgpe1ubXuxRLe/lgMRBrVHj+c4qlYlry89goX/apfDrcEvZ
14UInRJCH6Mhn3eNokZlaBpYdoLSicbJsO+8rwDGUfZW0RclB63ZRzMV4hqKbS2o7DGvDOh1Kzgb
iuxnt18ntExh8Shi+51u+tGgNRQjD1qrBJ5Xds7im+egqMg3xHA065jOgj8qnLbz9OwgpNg8blA5
wr+cdkYE0uXO7i/vXidrmRNoXiLTbEzT1qK5JB3+UUd80cP2mFi8YC+YWL7yQ4hTAk7dgxfurvd4
l322oV1zjONOP/sVWATL2SY9CRSF1GhdaoXGHkwV+n5s4TpvTwxMt3sKVRl0MtfLU7SXCdUEVkGe
QXDAY06bo1RhvnAEilCiPnf5Zgx+6hiKClwc+3IQKtsBV6LnNSmQYVit4moyHlPHHuBmJo1urOlf
skG0CZsBvLexnmo5x80Vs7KUmMg4nWHai9xL8B8APWQc+nGMRZExaPfR/AXXBmOeRVl6wQtc6Ujz
f8chIZYGi6ZCU6neLB1sfirsBswmXE6468uoOJjPEfux9UkX6bXQcLfrphTNYS0X66p8bvQUDHn8
+VqLVbU5GHU8H1Ai1MmHGrXbc2P07bRW56KHSX5NLm2uGUf2NZISktTkLnyffQeLecPZGJB8S0DK
cmExPABmvJrsas9m3xKL1oaEDl0RDHEuXneXq6U0zNuNP17yaPVGDDevNBuo6Gq5INKc/x2P4z2U
gMk+RC0OMV/YvJLjWLHjJ/1ROOv+qzu04snHh3pNW8mVDwapKENEOfzW9ejeXmVlolPpDpaJdgF0
aNyscYXC27knABo486+dqoQGoXLDnTV06DFWBWYJ1NMLMHygnshOmWT48EQ6782J+J+jFcce+tC0
X5/1gW3gDpjGD70FdtklTj1OQ9YBQ3PmNnBSxrqUzZFLGSMauzEaEdnLTMa+e3U9TXC2hc308DMo
jYl9yc0c99smRmi2/vRRi3SMxmRD3/4QWVVXY+tfI9k35NxUEfwb6EktwPpJZmjzYRdIJfMwgH9z
xM210nW0G8L8pt26EwPD4NEClqP7KWaFoCwR5g9XSlwbMGWN1qqSrzRcNtuxCS4lGR4l/JHoX8+O
ImIvYteF5SIZ4FYjzM3gu27ki+vuhI1MhgUSU33UEpBCki9icUojCCE72dcr2NVG15mGGbG0kLCQ
iDxgnzu5kGrTEp+r82fDdv7bH0XDvtOvgrRx37L2LBOtCqCFQmKT/Go7azIiwAuGw8JxbTEUhMOo
fEBBSIQNPSakjtF472pZucfCqkfvrV/7yG/lECgBlQTiPZTMCgjIJVqmAJSZB3utYQVv6SMyKEra
Q7C3htzW6lvNzAZpRJAvC6BbqpNwZaBBZqtJDai8wwjeXK1ktfaQFGKI7h8eF4GeiWmsnb50ShoE
lg3NDgeU15fdIOz31shR2O9J0XC77/mtNDwEH5vLzaFnNS1q+GAE/PK6efHMvBSDRB7a7zubHO7r
X/BGtVbagTzLxif/aO/CvlkiRRIelRKyxNmed7gxsTS9iXsEKnzE+WcY4B9bKkL1gNwN5i0kaoLP
+SYraM/6FU2MnOQBHzbPRNdZVRM7x4k4sjI8gfK46pBf5knU0j0svzSRp7f72QOwanWp7TrI+ZdJ
B/mtQdP3IrZoHzU+TgvdwDKTP5r9urPpKdwStbYtlLSJu+72NoMD5HG0E7eU+hqXldVZVrGAVmJh
wU3vA65iTNzVUTgHgGZNeb7P6GBZJduC9NYrKgqDM6ZSQZGusLI/439qZVsXz4NMhVdWTG9VCnY+
fsEg1iTpWTZWQlrVyPxomIuN60//M546+UQUMsmOefDotNdaDK0fo3xrJQUAuMpMastL/ui847Pz
7bwFDs1xaEPmpR/j1lFsj81jnZxaq3j54tfS2xL7in6FmWwftZ2NgyfH6RX3tTOMzK1reQPep98g
HpAIAzeG3Co5qJX/LRkm4HEsxSrSCYpsOvgonMvVjEMVWptFhIT+bN0i+/QCwX/PCXrG8crgfMLq
V+Wcr9Oly5ME5ivODHplZ87wj2oKlYwUzpcFKefYr0OpVbz6MP/xqEyqyc55hGh97eM5sYXgex07
vjwUB9431t0YEdFx3MCb+X54NT40JRGMZMbm9LAmnP3BVMlnhc98sEKhEPJgdp2g+5NEzA9mFW2z
UuKT/ZD3dUUKofcvlDT8wGUzVZzqg3O4W4UouemIWUcAOI0uGblMtByb3t3z/gpB1rUOcMYDAPRj
nzrnytScsqAA/wNxyOJN/ZUZZR9FR3EYGCW6rA9D6HKMQmS67eqx5WTBzZyPoDzzuCv2a+z0mHDf
A9L+1nt+E66FG7Pdm2YAVBcg+BTAaLFz0lTTNFnKs8aqng3kzL5WlDa6taucr3CQrzeLUVMX0Mmr
T3Dstw0FCDXap0jw7OihwZFzjjdhkt3qST+aX3qsWEYCGo6ZqWb1tMq66/fEQ/T1PyH2Z2xTi+6O
8wKwmSUenDZPUAggbU1a8sDqtU0wtQwjiDfNPzR9LtKRceRlIFpq3YaLHnn5ca93LmKOIgiqOakn
MR+Ksa4wO5kLGOx+poLSO0TqVxOZgJ0IlbL49I/nwll17rQ0is93QvkwEzhA084ssQh7MiidGI88
jp/noOhTJFr3mCtl17UcW3FC3MgbOGbJNN7erEAmPyM3t661nsW2nSuQLlWB2tSkP0p8CJPNHkyq
xbWWOJC07Zexfm7nx3R4grnu3Ss+83Ou+Xsxsv1wV+8iMK0JzrSXGll6b2FBzbBw9pP0QHTzqxKt
Q2A0G0VUzUvbeSuynQcOz4yr/YESsD4m21QFmQc/eYoRNZZGh8nNTZLeX1hdMyeLd11vowP3R+n1
OY5NzpUg2xfhmoNdy4yopGitc05SxPyC92brNbXo2yau8qXyDdjXeV930DyszMnpe0bVAGsiSTrA
g8/ACYtnNifXsbNy3e6PLzip634DN0qq+Fh/deVMmzXI+qJZ/9+bwS0m+IxRxVJQDXzwsgaN/VZ8
qV8pClb3gIHfA+GiXqG68L3H68Te5C7q5h1tp1/6RVr6XT92I5IyQaEmhrylUbL47k/tYO9I3yjI
HBR6bTvp8oJx3rCmBcyHF7pL5z8zBOMefaNYeQF/yHUVfEiolalrKAJKLp23vl3IiEQGFr5wl6zy
DWC0d1FOQrq3kqvF3fql9xBD77jOcRkl0U6VS73ERcZQdso60uaI0P5D548qrrBD88/Ze8wwlMWU
08LtVG9n9UsVi9E7LIqscDauIVXlMfP2wJqXirUaV5dbppxrEgKp+Q0uNDOACOU2mG2wpf3mcc7C
uYx2Adonm9UTxh38WNBoO0qeI9iUApSXASFK8THyRKEPZ1/KgHwGSxTy4PcYv1FQkYwAW6Izgg5s
TrslVUakVbyGfg8DJr4YJuf8YlLMcrTxGrADnwe94KezZLTkt41zZP8idvO+ZvSHGV++ZPQ1tF5k
rtJneGk6tsybPnnUBQTMt+oHuoOHPPWMyzIug7v5BGC7NmIezA31zFIpe8teIYe6zjNDtgHSL+mv
ghFVviZMVQvGmGrA1LdlX/ptegYQjb/w2yQpCiTfrBJMKtVllNI2VYxfkCdyrryWP6eIVtn8+kzx
MuEnHn3W4LP6v3cEzaDafQ24CKtXVSX1xICDFbyXi7RLBoUuT2nnFz+yJEk1M0/h6BfDysLPg1Aj
Cc1tdGnHLJDpf35AnRyqHF328N0NmRyNGSHpJw3dpEk0U/ES+hsYXVmnAEMCfaBltPhknNT/3CHH
3sG4Biwxx0nfE0yL3jGe03OXpJ+7pEj2WekyT9mXVi1tzLAWER14uvWGd6H0kPXSK1YonKvft2iY
u9bPVTwAPLtHwtvWK6Hfmrj1jZjC5mJqDLxjMwXvVUHM1hZuuy/aYXcha4ipmzIgyLAS1ItLTnS7
xuqgPvxjXkGjCkRRumcKjFarIAaqLQ2/Gri2wRBw6hahSajI4fdzIyXK0x+W0Ed44+0/AidRZDL/
WZzTqn2JSsSxWNLRHThWy56PGrdXnNccj1ARdIoHG2Vu4hjKlgv3lW7pdrZ2NuPZPwLoCF1bTc0A
VU/0eM2GwxYIxEPoU14giQdZxs1Zh0bpaHSYQrnOdXgQEasdQFsl2liU4ZYGtwv4+lvhm4KUXfgO
CkCsh9m8Tud6/Ujf28GdH+1u5+kKHXqnJIkvWjOTDLub5jV28i86fX5SY4IW6dptkojKHJiJlMOb
N4pebT9usex9e5BdfRy2taMFn+gI6Nh6FvFqmaDRRD2TAKY0hxCK0cX+xzzbqS/BH157pWdl+Mgz
8mMz/g+CpN3+XqYB5pIYsjd2PufncIb4titw+1drcHmnk+1nOJY16PakPnIULdAKccFVa9CK8Gbv
/FpHpBAzTbLw1Zz5tmBqo1rWER6KRbJBeUrYkC7e4sEL4QpjnYewKj0pj7unqeFS3XeJFWqsGzkr
C3E1FjMVnPs73aK61kTHQjeyEfBE+hTCpurWgkSr5AbDjoclxS59XihJBhxcx0lcNoxbpMCulJjp
GJLyaKeP3b4Uvn2jfHVTSeqkF5mWk4plU8swmCI8tMN45ZWetwNN7EvYjZTCUiSN0KgUrTybmZ3G
lvlzc3okvFDTBsWmRujNYU4eEXjYE8aoZyT5htthp83QsiYo6izr2O+Nv6Z2q7ahsPXbL/otBrXl
/C9+EBjnBVcQTnW7IkcmCBXU46xEtT7QfsK8MVPSoeKxrwuXM/1WhPn9EHsjYdDCIi+HXs+o250b
TR/4Y7RpZr8xiB1jIYhs3nC8PPN9jgzxqd/hu3W5UQPGRxoDD0Kmf7e4dtarAYQKSbsOBUloBRjF
nHIG1xY7RmAs8sLKkN3wYKtjVu3Zvva252V1PPoL6XZCfRW7i3MtGGw+DW+4rakxjEbHGR3uHEnZ
fbGq+JLyyG0HySq/imoiFUIVmml/kcPgoppl4ZSdDW0udr6UibuYuD8PggaMUIcdjpThxh7PAzJr
hFhwf85W3mX9cv/vz+qlazdLjgT0rl3skSpgct7cN6mn5isnBQe5hVNxBrKGw3EntMEibGUjked2
sKDjk4PicgPNQp4UPDdPFASaUozzmi9nFfHqnXSesbpBVDw/85nfr9UYVsiPmE6DCdBZIckDBgTI
B/Fm57F0vMft4ekifBA5FZbhI41PJiUOZ4eTJy5RrNNEsvbCgL3Gm3o8uhn/CvVyrDR4iLVXez7j
CfEF5njOoBa4hYEblE09ipfJaZRxSV52Mz9U8WxFaSL5gHM57V4cZOfGC3bOyshH8rnoRU28Fs77
YKwlEH06hhv3UZm3zGMXmeDsfCz7HKT7nutw8jkzDOR2it7Xu3XQkNSbGUcCKcRmab1/N3Z/iI9d
ym2jiccc3+Tkps2bGnq4sE929pss3BAB5q04TJxvtQd0nU7XXb8AnN1l8Av/jZNw0NFuMI8ynp+4
aPxxHW/G6qkf56JM4Fv5Jr4pmxRPe8Q6lFU8M7ZI+XSzy3krqL1reYxxZ69XLsOjgNJ+3BTMahRy
T8y7SvclUuXXiWzcCNfcCHaa4Y4fDoXE/TJ/9qbQ7Bp8FNKANniLGlLaneyYrhJo+PZZSzJKGbUl
GjLLh1NtchdYgXJgSuuHunTUG5RX9K8uOFz6VHpk//aDQ4t1TlNDIg6JddLAHGUrjd25GYgRarOc
izOMHbHwpcW29uOB6KqZl+zbpWkixSsvjLaFuRe/uwYNsGbdH9UIzhtUWu0vYpNDr0JNyM/CC8Hz
x2sNkCW0GExfvj5EAHMrcgcy05ZliNYUtveorndd/G9pHf7oBbOtsyHjy2lHNVC9Lie6zAQDHnFa
KFJO23q+/TogQBK1tTSUoGRSWGMXVPy8YGg89db7F3GsQRXNCWCKepQzSX0V3YRFUj4Dvzwn2PEQ
gSBbLkvbdArsAcSi1yr7fFL2PywzUTyehC70byNf2GvSyWgTiLxiIqo6GEhQ1byBhCmj960aZyzQ
N2WDHN49ZiAmjtNh1Y6IG86j3VrbxkV0D1ueTBOJv7ty/urC2DevC1y4RjkDjgFCH+2jIScQ+qTK
oB9xKClLc6BPCJVTREqbirl28FDzqH/E1a7unpHpHM7s2GOE4CceTkQm4hzYhewL5KAh05uuOKLO
tXGXM5o+oJFEP3RTtkG3SWs/Q3Da7HzuwPStVEM0f0RG9D6G0vZr8xQXT9zUbENwwAoVym661yTh
H+6HyoVN46QOGltCA8U/0SqonwJLZFCtqk+qR2Emq1E1or9Lr3DYHeqO1KpGaQj25tAYHDs4N2bq
S1woK7d+7ikwdjVNP5RgCxQpWnQ6ozS4KwU3anxhsA/Y52eeMPl5NukPrWLP6rDmOmUNTRhZ6huJ
qiHei3IdQZgKTHkAc/yL6HOcBhIRZP8Jh7US3T81aBKvgEq5/upkepTcDHSeurMFFEMfX7Atyv1l
C904CFyBizZyVg1pLsz9/kEmmfNDNK+p4huTpQGjb+9oggHOVwrH+dikhLqjI1E+7GCNeiDLtPi3
0/cMj9H9+osmQnJLiVyjpaj0N1JrhmTui8iytCmp0k+WtZSw/oPLcED8DyGSSR6Z+wds9+ZsFgY+
MLrX28xXi5lCL5qiQLC4o66fi8d+NFLhTDMNR+rCc6LO0TSVHjNcCZ3ytEQUJfTSIuz5FNDyG4Oc
t5szLvWqm3bGAG2CX6dKOUhe27v9zpw5pRQVpwImp/hni0Peg+dNOIiC4VPJ34ebc1CVCtuhI6Gj
FbKPlS+LnrPQwK/FKWJObKgsFoCtHsbirLXnjCce8uFlmeyn2QDpWDC26i33M9nrMdbm2pid2uGu
iJTcNxqveRAjPMTrMyFbvVxmLa+OhRE2JEu+mPw+bzwyBSQ21QRmQH5IqaY6mKsU03HQYyVmeeiy
8OkvSNeQFL823sPjWn2rIn05YNC3/CTIh/UKRyzna5HRvTUbWGPGf/YechCB3uF8az0OwsH3DGIX
lYpM3+ZRkjcYfueSciAMn4g+yr8qf7gE5kEqnjbvb6KEbvNcSSIKpsRd9N9q88WoOvrYQr9mkfTQ
UQkdmo0PeC4BQ/1aKIBPVDpK5rfDVytFwbBmrAKoMG1ZjvdOpp9LioJMtlkfuh0ba4vk0yTEa7vo
L16HtsjRYOWNJvEYYVMwJHgl6IafB2bHzUbNUUj4tHvXVBgYN76fVhhwEqBwoDkl+WxjkWU+zFiT
IyZrihIf0PMZkbxMcWjts+lhlgy6DjJRhu9CS8qk8u9Co4jyAZ6LVOhdbBQy0nd0VfLtO8+TJg+0
NAU2HmJDNF/gPLBUBLmDU0wJiz1e/DEQgZlTZGf3gq8B2WfP/WtL+5AoTOAKhGAWUiy5S8Or86O6
ZUD2PPqf8eaaQAoF9uheuxfRO2QpNK11G0YZCTVJ3RouJdjZo7gY66oqYBPp04jkpqZI3RZsV5OB
eIih+1jsO+R/DZH+8mveIPj2FCMWdUTlBJ5+qq8pmDHQRKab2/HRtyRnH2OsPjS08RIdOM61630D
6qvWQEHgh2MkU9EX55rqV/qWHdrjK+wsF7mU8A82qHHZ+l5zBSNFCLPJ0oLNna2wkqoeApOyR1aL
4pp4kf60FYIaEoXa6xKaKeh0RfGxBVUs/PZcN9+8nAb/lF5ebW3R6+oTsrX25eCtgfFi6Jm8ECIJ
7ntZQ3BLb+igL086/aOgrdAZu0xa9lA37dHF7nrDKu1BQC4lJWQvI2/5XOgQrSQdzNcp67mRqf4e
NRxcHnDSHIpwBL3Oy7HMeJt2oobb8icCaPDYs8ERN+sIf/x1d4h7u7/b0PtPsy9TgLb2PrvZ7Dg6
4DVXr7AXKJp52th0FDuZPrH8jgMTNrPqi/gm4mbryty1B0BG279eN7fUxy2VxPb4Dh+hAgH5D0a8
6F+x3fwyfjyMSN803IM1ZwRr7xHnZjBMJY2uUUdzKSa2hyCIf/MoJURNRts/mX4qDeYXoPSap/wL
gKCeUH+vq8Tqp2hih7O6BauVRHwAmb5edLw162F3pJdFboN8qRvw2WfjGXUoV2p7C4pjyTT/kFIJ
7QDauuMujcsTFOHnFiDv+BZ8a67+uecuH+7HRbwyVgLdcDy1p0etxA//rLY64KA5x/MacFrnQTWE
6TDqjOynAk8F6Rv0uYM5wziyqVOure3dmkleUUvo/+Evm6GGZ9OFGGCWSBTukG2pP0AOCKOw0XTF
xYiMqTB9agzrJ0aOhHXmCwxOwR/6ypp7/OkwbN/TAw8c2kvBU9QxUjpu7dS6xKyHVMBHfvTeVTa4
4AkZRFOpsx8bXrq3vhW++EKcOyFfdMliQ0R14oUuaadBUOdr82WVgc5rVR4wlXXEkq1+6BfhAWu5
MhN0kn/HuXjQ7WEtY0uDlYU6M/Aw/3eHJopl6T4+FJkDnQROWwqqbnRATn8BjqOrZO9O4m34Mw4Y
AOR09WpgXFc3LFZ2xGl0tLB9MCoPGFk+UbtlPNbiOu4pxr/AfkaiGSKPbV61rx5hSJ4ROFRYgnCW
yCVweY7Z0DK1RqxlIDnnMHblhs2JeynYyKMMdhRYszbHVi3Ir4DsQvZ4O9wZXRRqMsi7RN27EFm+
yLDtaqQ5EDsQCx60/+uHZRrzn4mFmYB7ZBYso3zYRx6V7moyOt+kE/qrKYiayszacxdX/PNJNk/e
n/Ni3my+oZg6+Qe5BEY54jcrlI06VChN9XKojcg9m8cPIEJtPpTioU7Lmy4p6njppliaw7dOpDBa
tUVcrcNyy5nnKqK1YOmhQgtVRZ4cCR94t79GnRIPCRBXnyQJ6051K1bbKKCYA5gQ5CCGFBofwTz8
5q3XtF+yQ8YRV2/SO0thQdzq+UUDVVTDM5M/EQQxZl7FStW0xQbiqe4g6N53K57WKIT+025011kb
k8UReLavVYd5YV2QezyKRkrvcteYH5nDE4a5d966XGymXhuvuLcNXnJCOUfAdDDjrxmtafEf4kIQ
HEoFIX1QVxPrW7f6aWGsnE2tdDhEBxKNn5hRk+fckhe0JBc5LOEo11hF4n1VdPFMQqY2PlGnGmFW
6XhzAe51ylVV8M8cQnKB+geEUPw3BmjUoOm+SNF/N4Dg82M9F4UUK0r8Fv37FfjjrVWMl/Jb5que
cocq6wO7e7/UY500y8IZxlxf+ZTTVXI5nWO+sJHQYaI/FjfMLPnHQCffpjcq2ZcoNyjH4iVsXGGI
ccfQxFdaZkdXrITk3O81iS0GsenrYw5I6TaW3VRjCS3HUNGesjOjLt/lwTkDedj7ky179A+oyhbf
tHEZcx7UtueUSgSANWxAyl7SKpPFsJuxkESnqHYAwFQl+NBxiDGQS2Q49wAVjaYhCB//5pIQfku2
eRLV2A9LM+HO7kqcd6JxvnZLKLGn05tpjGNyo/TJvMkaoo1vOgPHNbs52+W34eA9NEl2w0eT8b5i
/7gpags0B7M2lI0NfeXwoV85IiosHVpVbe9k1XJXRMmoBRjoAAiaDILgLAlCfYKKTUOLCXLTgQfW
sRV/gTNSBqYg71+hUli3fyr4BBip0zpAZBGyCoPxWu75eyWbcfCjDNl5cEzvbyoc5FupBjAL0fuC
PC1sZX9ZoCEpu4PihsNN/PAJn69RJTM7IFOFqSgZenKaJvDfWqBJdo0VzFLvZJAcvmVvDkOVK+H9
t29gzfoSJ3kVnZZBPKhz8QbCvuLqQejcUJHgKgvbDzsiQfOm39sRVottq0peD6WvSzGcrgWfXaxA
CmZNtQ0/D9HV+OQD/Ui1kDycJFedXJKsGS3hR+BXXrZ4ukdiNT+6AAt2Swb1wn2F1y7bmRkxKDCP
jycguAjUb2bUkzAF6MRFVGed44L66D5JPlMrwCCsgfxcbYsAV2VCFpYgROrLbLTPedy+C9+z5phD
BYj+gVYzQjP20CXkw6c4wOLF6axQVnr/RuEKk6yZbgCRseiLdNosNT+rlHZ7s17d5x9vjoSl9HWH
26l62ee3Ts+YI72muK44T7FeF/ruXGjqDOwQhxMfBZU2cD4zHMHl4f7Q3+CcZY3/L7/ovPDp5B7q
cD00QvZdM/vk01ICIfAfpHvoSSe67gEtWsRngi7wQWQh5OCHyJkbAX6ZfjwqyJgDz9awK67eMhwR
xOgBsLBEC5AUyUhtS/7p6OxAsw4DLf46akdhxlAf3cZ3xmixWgVv0532ZE6ErCNtw3GHODYBcFca
YL1B2Ni8HwJOT8qMDzkElzA0aOR7u2qgmMKVo/2vHv2ZKY4rjaUlHFgMx44INnIPFBuOSMVnaTuw
ZRn7kBY/KAxrVmSvgGiS+OFcyfvrhfizEKexZHeEUa7bnqz5ixRB288xSI4+gbZD2aIZ6BKm7mjl
1iJlij1jOtD+ZQeTiosUyHmGxuQSBmRPeewQuqebOMrN3hZgi5QeUHTzELDcSsDSQHxeEdj8oEVE
Y0ZyaM9wImt9lbonH3PNReqDeQQ/VEAILsrHZKVGq3fovqp8dbxF3bpsoEu4sqfT0Qyk7cFtRsv0
LJi3UycPQ+BcQ4Wgo123WH8hWay9bdi9rM0wHXYfKod0ahFyMfINMfcw31T8pmfWjenLXCSOSw02
xkkuOcx+QmBoo/1XQZXQphnxkQMny75tI0oEBfLpgV0ZksVdLuQ4u66HekVYrnKfc/pP8Cjgwlci
j9spHu79OoCNTp0mQAYk+B/S6rVAgdrt7ORpPsibz+LFalE6wRN4ELAYmBH4CErJHljeo2avAt2y
/lEAxZ5psKZCGxPrqCx7RSx8f+eNWCWG4bZdi+9td1lycxqIrgQth2EXixMPsvqnXz0AG/ufp0SS
3NAynXpxIG3fpacMrcCyWbgTajkdXlw8usIqabPZdcidBFNr++Za/jYHtzWmB2d9JzWQXjSkhPj4
EJ90Jig5iivVUrJhsSGOjxTUZm2mvrws2R455OT5jqVLWCR4Pkf2JLX37UP7D/YaGvKrdjyFXDtx
vlsGMmBi8Z93WT8FJblNriUxLHOzY//wY18dooh6zgfMNt1xDGeBb7xoE5cYM6Q9Hmav45C/pO+A
d2Lvo6/pk4pWRpLGUpW5DkY20k87OKHU4AstQH+83aDy9ZzpmyqoRKbdSs2br2sAY5+A9Z/LmgQx
v+Hk7r8hbe+WAWfRkPZcVBJVE3t+01RRoY764SvuPNihWQ1VYxrqVZlLnnCRI2zOh2oM4sdvRjRv
1zbXqpLbkKrXx4HknzFoM9oBss2C7PC5DP5u319c0mhXkqSNSRhiQ/V84bk/sAI4y54ol27VMbqE
mwZI1rn66JI59T5QGEOe9ErNHcFsU10EXdDogLhpj9fn7wQe9YXLaP6qzMUPRHhsXlGhcqRFqVzh
NB9yRz4RV6NPeH4kEzveBRaDu1hEW2/x1Mq9SAOuw0dn6kjziTaJhbkTLRnp+8VBjrR/owSms1Of
f/msNitYG/Xh8ZoSpCQthaC58wDb4dR8lQ6vdR4vw//hbw9ecXLFUPAimVNEejOFNEZEYQYmE19V
iQjUsUhi9IfpqbLqV/sPUhC3CZXZASKJa1a35zAFqMnqSAFkc3o89MFq2+0ex5s1oT/EabkAx/yh
I/9qLS+8rZsMN2nESLoCdr6PF9bkLJz+dI+PYbtrRuc9JtBwowQoJ890Rej/egoBAsoeAF+l7e3w
+8y/XG27bC/G1Du3vKgqXB+R5wiw6QBZDz3HYTYCVdsPszqw7tTJmQTUoCOjSLgKfJJyRLGPf+Pw
PXOGdLTzilIN9SFHwMyXc+jypc/ZcViWC1LKnq4o8MmA8Ss8VkGKVH9/9dniQNCUVKxdb4Ik144s
6Se7Oim9vsF+R5q71dSHiZOnXJLNgWvawOt55lmMVifk/B4CT9txXx4G4xzYS+EujcqS/3iO3VC4
zxuj20FcOQQgLKYYpnJo1qU2FRIUtGECnFe3YszNIH57diGEU6GzMaW53CADFa0U3xl9Rn6+jFeL
txb7nzAEYXWraqbI7iPRjzwjJsBCSruxAhMN5XEPGdQsTpbxIxzuuCV1BVSF0pp8QYyuRSadQ8e8
4Mx+3Cc+/sSECJC+9rvnp3VJNY/RFmGwSeYhH5f8+/1Jz17yiK+Lc/pW3iQ5+Va7Wim9FpcD2rz1
bJjApe16ZnRs3azlmjrFmSX0A6pQuVeVw6f4dMtsjZtxGIP/DIAhhvjZg/H/izWyRXBPHSXcyphr
sT7pXYuQEUbWYpKlgADPjXNmCfo9EV04cjItgD8w9S5eLptnpOB6GDokXoDCYQSjNK2wOUbL+3zz
Av0JRnLUmay5iimAIKy9uD3lpRyaoKPGMRWcxL2U8v4oLvnZEfXIqN3zICVu8cggRb2e5Y4zB/hJ
jMNEHzHOkWAzoFojkl7HtbIQMeaQal1QAfLtvFw31UVuiohNnjTRhf3QM3iNXESsI+IZI9FAyQlg
GAaxl6edrN9Z1jAH34H8AAcw3aYVGLB1XOAptxAY3a3Yv0sKN9plVJqQ/YzO9I5CBnSonJFODLDz
j47fajwpbnaJVgiHSY/K8bKGclTR/bDhLp7/rOUOS2OFPlWCY6a3nIGQfUICgweNXp4K4I6sGoU8
737jo6RoFqToIyzWtZt1PS8lfuSsbE32txcYJQH9NFm+OV1/CdmU5di5gFhBAOvDc4tYng2Xe75n
I6goxI29z7jmoJTzppTMjNo8T2pnosTsPBrBUD1RHUgLH8ateGHfxjiYesx1lKkAz5KeJyy7ZJpq
jOZtJoiNcofOSS10TNYDqKGUmSMpWwJBu/iqOywRUpMPmKwu00GyHJ4FazY5x7cuIq0W8vHoIPI6
n9phwF9+17En0j/GVlad/h9wN3pZ3tnHZODyF9x+UCmlxvO+KkOqzNdC8V6/Al90Rqj4ByWxt1bk
s2/oXuUeaMD2a0ta5+gOBmsh0CVH2uEUeDofTyvWGt2erEBoFod41fynIe8D6/R6En/7ZUw9iMPY
P1LXAIUudLIvZ/Oh/yF3J1G1F4T7CFk68cRJa3wZ+yKd7rsM/Sssief4lxRsypQecS9AzHhqUhms
y5XH8Dat1RwlVqGn+EpvBHxNw9KDARHYTDgjF9tn9Autt1Nu4hRk3WOxq80DhA0iWjZ3LZDSe8ig
e094s9lVAWGRh6eDCtHxQ1jttYH2XZGvL3II5lFsGzGmNbdvECYZ6sgoiJdmNDUXy2TVu7IPJ8rN
+YL2G3wQHysl/TUCbRabMjOkO9om9iPBQxtQnCjDbzJoveddjkN0+HQMmy4puy2nHwHjR8PF61Tu
YEUhhsHlx8M1KHBysGEP2JmS1yL0SH+a27PYmpnv/ysxRjOajC5ecbFXG10HKhKhCCVg1Kp8vbcK
pFJinch1lc1vGTPUnfEmDYCtfm7Xy78LSgd/rL6sLfAHsnOVpOwBzNqYO98GHQA72FGWoCpaliqu
gzYj06et924FB27Y/T/zGOZf0ZbSUn/y6P7plZ6RvZEOnhyrvmWPZ4kH3Hov7pr4A5WqY30+B1Q3
g6zvHQp49bF+n4pQk7zIRYLqEwsOe1IZU8xD9U3QDGY+QMN7BySVRmsBNkkFfwPPeX3j353ddTay
Rof0EYPcO7zxKxznxPYueQQOf7V2xhHdiFBAllRopBUh7Rim8lQQjmGx9s9jIfQBkouQQjxqYj92
i5By1Giko6w93u6tTTanxtIT5L+oz4/hio+2REvJDjBTMl1ka1U7AtZ+r+L7PO/IXR01wgeaQL+G
BkIMqZdxsHSnKOaXa9X737Cyh9aA4nm76zCEmA+a1w7aotpQh9ciqpJ1KXqGLZ1T87PCmYwKPtaO
enWgOkCVRhcfzx4K/NtkrKN4RdcHQGBdM2l032lb6b30xlUR8w07FTngxTH9AN6ffvQeeBTJbOWj
UrfEIlN7QzJicuQ/bhL9rOw5Jl6NxRvgMe+YqxUizU1Yaw+CcPTW7I+hnK3qFlt6LcaQozLq+yqR
XyVmQURyTobsIZKsytTW5B3fqouSu4zqUcppmn26R7yGUOo13QjuhD/YGUNU9juemFJMSLJWe3Yw
L/vWULgJo75I+8WaGeZ7rMDC6ee2fJNtwe3zd/3NAo49oJcfm+VYIhYIerFgX8MUrvYZCOjMBDhg
Tmpg81MoBD+yBwoA2mqhpcYSuoXwBtd34zgz0ooO6kz3iS/SaUxtViPOx31ua28bCHiSfI6fRy12
1fIBvzX1tf+Gawr6k6X1rtreZVmJJ5+BroOnVUJDTH+7zi6rj+igzerQcef2zNkQxtPStvr8gU0l
AY5QQfaZeXpA6T1q/w/zmA/rnq5i/3WHuD/nhqqCkLHyw851WgIUwhCXT2D2rV+plNwlOASa0/AO
rBLMbZFD+BX5tZ8PKFo0Sy2NUeW+YffYUWD7v6fU+vlC5DbwC+a4LWkc/ijHLl/p4A0VCT7iwlVN
Bk/K+AT7ZrfGJOcQbS+XgnKCs7zjErcPQqlT85h2hVLCbkv9CYCMw3CRqfi3jRiAOxd6EuB8fcqS
EKDAtPMn+TpLxiSkwo941bD9als12K6zT16E/Ow/nbw1DcMPisTAv9VMY5I+IL7wONKjQ5qAKMQI
FCNGr7h3GYGhnZRgj03srDHXd8IhdKfGMH0Oxpp9jaQx4jmHJ4LtLJ+/rVR4X0MtNBvPONgvLeMd
g2qgAZ/XJzVL2GUWd1CtL82Wu7urR275uNIwH6ocWUNO/4gOEmkh6OyQmCkGuUBgwOz3sV8qciXi
G+MHF9FXXxjLfnsGUla3jj7mTrVim8ZcLqgW/lo/FSIdcLQgf7u4vv6/+pBTXNox6WpKhwo9clzb
oJWPFqDs1+/sjERd2TZQzgb2q/IoGCAcqbgV0SltmH/RJ1buXfgsc7sEuNDIlYacxagectBce/Vf
Y0PhU/x/UvyA2GLJF3nEY/GVqqcpbaDjysTXPLqt/wicSbmSDmGeWq7iHtzXiXf1ZnxyqMhn3Qez
laI9+3U8jww8scKVX2dVE1OC0RNOSaPmkcI7lygJMFoQqjsEc3CR3KG1iova6tX/mK1dPwx148WG
Y2EraKcxmHyiL9TRtimuVY5/SbmwsgLJJP3Cupmk3V4F8REHjJK0nNgFNOYHqaeEWNniQx0xtYWL
Czp4D+uhCyZ/qZ+sN8liwU9mbQSSZtedWjI2CRtmn2WFc1uDUppcXXQvI5GsUXfmilLfmh65HSIx
rsTVWEq0RpVOxSm+ewdhG1hfoChrFIQMNkHmm/kyrSMq2PEk41qqblmfTIucH3YQhScozNdi0Y6u
56DPR4cxcYe8dsu4jgYar3ogMWQMrayUZ5XBP1YkfbVGn1rp42EmjN+5Yn8FMV9lU8HKRgHbGkZi
O97XhhPBNzZ9txAxqERKHzU7gKl06Kco06o91BAWlN6wYQ+907Pxk4pFOqBLcN8I6cGk2nod4p3L
PaurXsWxRuu+c9hRYhqxOFNNzZBzONLSg5mvDSsSBYIiLbOSd0UFnu8Cj+Xwow5l/w2dnCSAfZGk
srNtoWXmNrgVnV+zJ/hliXUMmDLWz/FJ7I/qw8FYX24l/2hOdOS29woRhwKDg8dCA50EhtXQsoQJ
jGgsAA4/lyTgnv2IQNb6VJDeMRA55+T1/LJVHrbt2bFZiKx33wkN9eY67Z/GgerkaN2fM+ZTZcxW
Xq0bta90UzfJDRiFPVENV1Kzd2QQrA9eeV7/ltApTKxmcvf2fZwPcPzzLyREv3NQ1vzvECAgZWe7
7sZOgR3E0Gx0vrvBseDobogfhsVAQuymhYOW9/zNFWSHW/DGh/WyhysKyQ4dHYnnh5JLnm4gDxf6
AIVSq4n0veL0tusgb81pp5rOeCl8M1BcIa82moACKCoszltc9WXag4GGBZfEXdm2Zf1UD61cbRdF
i/KTxy8Obc/dFHcojMoLRq481g4KW4j5mqXRWeLKOSeTCvQOzSKadK7RgP9PXOqflNC9eYCx4aFj
WpOah911kIBtJp/LghGMDmqBdpAURh0qb2v9+OoTM7/iVhslPLy17EJUFhrouV2yPPbtQdaPaENn
Re84ALq8aSc1Y0vy48cViHO9UjTdXRa9Q15LcRtwUnjrPL9+ccls+dmdUBX3B2EOY+o3bQcv/ub3
FjjMfdcf5ILDdDUU9L6iKBYtxGkkvy0pMowAJJW64+gtLjrejuJEIkn7IBJiCuWXIRJM+xaWy2I9
4xAeb4VRWaswp9WrR4zz7HaS3EU6HZf5/kdXbdTOjhk4UQYLWYyYiNClC2j18CRNe78X4zPmccoZ
2oxUT7V4i/hkGzfY7b/uURPcjcU/rpCZ4gpcjkI1cZOZwcU+8ZQBl0wO0/J9f8/RJMKME1Kw2XmI
ikCX8a20i4VFL8ZX70TDiGb2xtMYqmiERW+piPHx3I6sHbiMeegX4SNB/mSn7w+sjP1dXrT6Ax0q
Uz7DWL/hJGwHZTszPUbiIik4/kUTtrQHtJG2uO9PDcdFfLs9zNWbeoIeYqnHxH8Q7KZbsV8yRO7S
q5IT7qjOaqOqUJNgPFARKD/DuFe2WfbgoSPNhMoXrw5BErxoLWv2leZVjRW5IG24woY9IGgGlo1s
F9ueHzhPUEwVcZsPUvSDu9cXOo4QwLLfr5eWn5qnvYi1NFFCZcbV1rUvDL+WBhWSmf3mSRHvlLRV
mxsJiuRYLZc3a5h13HiczFnv0cqKgYO3aHp5/hV0aflnteemkoUtfF92h4GbMEplnaUXBFDZ9mjP
J5+zUdiJGHEWCIoEikZvnseiPlLYGmN+cg2rDZJ3KZEnqzHVnSic9/cP4O4Ec8vmX/AOnDtznqND
rwAOJPeaC5HbI/izx8t3AklfEM7G6IuFWZth9tClMa1RfJzEUUOsUYS4TTfKh8+xpvZlDh0VKrpx
ijro6DUMTv8/RvyJMjaYIB0hoV0Pxw1nUiuD4xeSdcG/BF9izfGOIJHb8kaHbeo41slQRXSg853X
NZO6ZbGlv8NwIJtkQhxB81s53eWMUiAhJZy4Za3UjH/8h3ssjHpg3XPScC0GMV8SXjJJjlpibgPp
klYH5jsaN40/IVC6gwbfoqyOn7XLc7TrPNCOp2xt4nvjWI5SO0LT4dWCsTCBJEKBj2sC0CTDUk0s
bROjFCXp8ApZOtgw/YR/dZqQDGQj6ehPRK+ogZN4U5mwmyyUDCu5dAWg4go9SUjIB1kL8TwawSGp
mfVKuYERYpsS9NmPd6xfE3wLwl9adCP14c0VkR8ZcHTYLLB5tJ8urmdRUdwSIBCzRl6azPQbLjkD
tDtPGsw8dq73vbcbrBvvtWl2TYpWMmsmcUXphRv0NJJm45MOppKBD3w4PLOIcYQUQVOUHNQNesGn
Aj1fz9Xe0/GqlHSqJZp+2WCpFGqxkOvoEwEBDJbdmUt3zF4aArfgIXy001nVi2e1Uf2mzwlXZVd1
UB5Pe5drk5fRAsZRQu8heK6W3Bt5kysBJqEblduYbgTCzdKYfIHpaJxNsWo2Ah9Ngub3YSfACW00
HiwDiot81XDPEuBBTXmP5aBhNK/PTS6F2ZxDV7cJXkO1ZOI518pSTifJNeGP5sMKCPA0FU8oy5Fl
1C7MPazK74IH1QwKW5Pysm5RUzKFnXqW/00/CvszdUSOKbhm3lLwgFlTJJLiu3s+1m+8hRqD1PYd
17KY0JjLp5TW68QbBKUlGvPvxHY74cy6w2ySYuyaP1W+js0haoxUPaXlDlt8nIuASH2e81BPElNp
rS6sCoP63OYIif2jXcdiVwaBy4btc0s0z6A83el7kcqKahfcqyzZQtcvfG/w8Sa+0zUUtinkuPUi
Llu5e+gupu5y9Rq7w/hWBtkmpKzQklO5ielz6kDHUjYSGISL/niaI4EHIkzphdpxvodJ08jMQLGO
FMqKViQVYtVV15H1sIgdEYo8EKuuozs9A2V6at3NGtYZ3UKaaamCO5kkaFsK5ndUyUA21N7CFewc
lLdbUiSFQ/4KakVJCo3eYRqbIdM03vuWYbsPdkHhrre6KvInok9Q74nxoSqPC+VULjEp9D2CjusN
K4I4iXi0klNnobfI8a7tlSqJGRYn3NFxB6lqvnfO5Toiu7pXokZz3UVUlzxLJQomuYhuDC8+yBWW
y/7WmM3MvNdAaloJWUkDzTjff+jEWYRCvuwO8IEQbcnGU9u/i4upHcyW0JjX18Ad9GwUzK1fPgyc
jvNRiWvJuSQuL9zzJScaUavy3j4iIZiNoHBYambg1ljZhxQLY2Lc82RyyO8JfurVri+8Wuy9X291
7dVNVVBmUkv4G7f0aSOhnY2QRl6DFAafouJ0XgcUOP7XgCwr2XEX5Cw1Brpcn6ap7zEaIaFOAnJk
O+owQcs+ZYT++kwLjRhjaEInenRYVquygK5fdRiTjx5j7C5TJhcdGR/5hCzhyPsFMHr44FTw7FD4
eYGBrFCZJ11ixDIVY3tgZLlTAnpO0H0MGYbXn7gQg6OL/E7IGORhXwcb+73jZhXrHshBlpOaqTXX
gK/rNz03WYsw7Jfjt8t/dYA16elWZv0V6j9rATdA6UFSuMTIz+efCya+8okrDwWbgD1nFBmC9pCL
ATBc+mBpD4vGtsyoAcjOw4myz7aL4m8Dg2YE/5d0iQ3QAeurMC9U+3gCG4LYMibuG7z8xnTbNEOH
949T33Qwd0L9/dI1dqb/FCIRi+v29R4iN2AmKfvp9RfE/yVBvGKGq7NzbNoQrARUj7daRF8rVx37
khFzFtP0qUJ0hGsaX15e/r2XggXAEbPKAqG8hHSyRaPwJeLs1lBfvTiBfWxJlsdr2motNr83HG1t
feVkT2hNp86x42fh8noNyhcvnKXVMe6Bl+XZdbbrT+tBKokeKr0P86ezjHi7MB9XAmptstfdqqDj
hmhCxPZ9z/UNqx3sIGvfaJSpIJwjkJoBxUdgQF6CgUoH3VIaTf9i4ctriObtRoKhZTgSTIakEJCt
u2hwn2/Mtm8KlQRb+LxTZAiNXC4+hKmWRY69fYQGjJU+NCnUcCTCEwGbIJE1hsA=
`protect end_protected
