-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
oZs2Li+F9W2dyvAa4xeFmR8KeJps7SMEdsmbvLl1xbZvvNRUAWkv/ea/yMctCt8FQAHs1YW+2Ope
vyQoE3OjdOBkwZC5ErzISpOZM4WWo9u/ftRXFXIIopyz+wq27uZ8WlIX4urpdNHYZ89s7XQQjpfA
+ieaGEZAQPw+qnmbpZJo1+Hxl5YkkGmvFhRyMLZznu5AFlUM01FRZ7ln//2RDKDFqNFxRzfuWqXp
aBmNl4yT8xddbdBAg0JH9e+vrFtzDXWrjkaRdq1rFEdhflZIuUTrbZAFEJbltiQCTx8J4/yOAq3P
RINLVRqVozaCQU2GKKSJkEkr51M+k/P/jOAFyw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24704)
`protect data_block
C9vn3e/artufuk3SzW7hUz2/O+f9mz3ZPHCE5Eag+ACW6cGn3TyxoxZPfPtU44gzggP6I4MVRZ+5
V8glja7o4HdPMFeVwfVTFhF5EY3YWpqLeCMNTYAAOTcNCDf2pfm5FazEPj4PLFNEoJ3YFEP9kiUA
v4Fn6g/BvxfpvwaERVfzhf/jQ7qwsz3/pTLLhCR6tEJEIzSophSTJ5bN5FWiCGrTI4VUxs9EN+oC
hTuTD/dD1IFzLF5y2yomaVwygVXZhNQFfDdDpL4rAt+mDodWpbHdv0FPcNkwP0nhOfmIjgOkpDKt
U1crhP2rYY755irg1Gk3w+QZzSrQm5WGo8wfRfxSrPSYYnf0nZFWUTGzmfZyvkTPhwv5MN+RutB4
4IRTmR6pHYmeiRv/Ioe4fdL7SU7YqzJyg17HYap9aayFcCrwQlheeCSMBaBxvHL0//FTcL5MtDTz
80R+Y9sZYCj3OoXtOESX5Znkc93zVtGpZGJM9xJUWRrqhHdrqUyJjE2j1M8aQuz28RCxpS8Fbtbb
WAYVjqkPH/JdDc2fc/S2eFkCu4fJZwmQNc0sDfcDGiN35DbxF/0DrFTT5bsF7cjRVawZMQgDp9OC
P3XR8786hy2iu4apzy7uYOn2esp4un0inPy/nwU2DQmNSLDN9Tvwq5z+9x3IOZahVCdxVpldWhYv
lVGLmTwQNvCZ0GQeVbDzswQsULNjNaLDni+abYgsu6JbQFPem9RUwdEQ3EtM4s0vxwHCbD0XfYHM
sNWAmu1XV4KxBQRkhve2RVcTQc41Z/xYR3vSwG04C7TaL0xFLqSeeodA6PYdWdNm9FAXqoSgbeXA
0ddoM2bSdsPRcWQ2bN0PcIAww4hUqZI2o5wEFg5aTkfSVFxS36r0GJmiWaiRtzE+59XZm7JKTtbJ
CEvI24rduTkN5nDZej5RoY9WiBQhGPU+MmZJK2z4qvqdZUI9yjTWoThZNd514WeWftHRGF7pMK3F
CWaq8Z0rupfMSkmkJyYmMlHDE96tg6MFA5kuh7CN5mgNBAhgGkvOZo6+7mEbqVSvRnc8EQTFIyUW
z027Oo2eJ7LO0PGeSeMPR8JfvGoNwaJYwNqqahqicatqP1ImAR2WvL25vcNAHwM+1zPzeJodvcBA
oYHwOWCviEfMiwa++3rIUrHP+XVY962GH53qg1aL8khoSVdqUrSrkk+Vh42Ww/sZfzIG4o3N/zEt
1JsVxEgqiYQUhtNqzjnPNJqivi0yEDwbW+hbzH+dYI9lN0ysoeyZsgI/ehkQuLECuJXA2haL+zWT
OBQJRSoTW2BJF6cGbMzJVL83kjRuBJ0J79IZOa9900zD8pn5/IhKU3dMFc6qgO8H0b4qV7wutbw9
JpPCb6sOlWjAxCofLtjsk0v1Xxbr/VBTME5/4c1ED3YwdEON/W6l4MCucT8KzNny/G9jG8x3BvLg
svutTpl4RtY86Ueko+3d3tbJKxpFLmzVY2xBb1c8IADyA8PZETyEjt8smfF77V1rLraF6q+hbW8o
DEO7ZF6rqMU60LZnjbo5Ir64ulP1q/ZHw3m/gEWD0A5zEJjN5GwswuQaklqi61hk4gZMJQ1XbyJ0
bEX2IScyXYL+8X11KdM97EmFD6dWVPaCoEBFfF1xoltS9FZD1sPNoAZh8atyRAOM7glHMjUrjkm6
i2idj25jBop7N3Bzvaah4oPSEvfzcNkb9oVH4TKe9etzz963xYstcnB2FUsIROpGkkgkjn1TM3pE
LR4ofm+0enr2ptEZI1KocMH8Ndfi3bogcVMuqWGFTFuk0t1h6bjRUSFMY/vVa60Bu2QG8iqcLRFj
fZ76w5seeT/pJ/tvCEy7riTJLdcY2mdWSTdAsA98zKuNNO5UJW24AYhR0RCKrndPTvtXa8XYukra
YylSk1wHfKw0X7w80WPN0t7rOMIDthTuoyoyQ/BCusJUY5TXK/x3f4s/vyd/CFQeJMLSvC20stxh
GeQNWJHM23Uk7ZiGsBypPnVeCytW5Gx2atKqln3D/UbK3Qriz3gSUOJdweebUkyUwBcKnNRQZdI1
IZxJSSUmA2h/edkBbwgk8YxAWVHCeTEElYGpcVVxfSSs0HLW8zWaVcoRYTG21rjvxD0r3gcxRIZr
0b4DNre+UYHAGZBE43/cJYeZiX8XZV1Tlk1M9WSrTQGqKrn2KAiIEE9W3RXvwPwwBbopPz+NpONR
gmZwv0nltphraau2gXp73m/q6G2JY8Ar4xBur3jWlP3FBiBOTfJOxl4XaWAzIcHqvn3mwJ91QRCG
mJ5QwPmGmD9/3Q0dugBXEuYdr1Omho1QK3EOzcraNOg57lwZEv36cWgbXKOwqTvWYHfMBbRFkRqD
kJgpC+d4WiZqvXumRwXHAjg13Xjysz50IrM8OWN1OzHi4c0Lf8I/PopY16JKeoojCEDuCcLOjZbY
yFiOvfNPzCfe9sukNmbrfGJPDu6c6Iw2mEfiMVAXPJRfH7klZwcwqT3WQ5kk0vwrb7J4YIjpHE4i
zyDOVkad61KL0WYuHCeDyoWSqwEXG6/7lFJGqO1h9nqakDUymI3aLpCtc6OKT1m6VSnBabwgbUDg
qWI32EOJcNKpX6uYt4SdVTGaJatvF7h0TE3gZmW/kGuKrvDmZ9mkb3qALEdDXuGKb6P/wbuWO95Z
Wb2X7BaDzLJFHi3vFSeCrKvqqH845us+Yw8vBhppmvL+Ysmxa1B2tiXl/jH+4OOXpcq40MwjlyaG
WGOaKrGQkf6oRyE+KP+dqMEuE4XL+2gEVp58CoRg/ttJCZgMul+sc+UEN3GuPf8hP1MHggvCIE0A
wMUJUgKKBKPfvPT0Ez92GXs6oDzqVoGKjXytW3QCnBMdRlnYvHUzVSyI/J2q5B/xaBEls16IfTbq
rEvH6MqZjAGogbr1Acl1A6LuYes+rpHFScIxwrcEdeo0VQV1SXX0DortZmH2UDiME8gYqmNazC9H
G/Ru4DvQPxTHt4mwgFO+X0EoBmHj7xFKnm2KRIoHEQD01f+ZScAUu25KzYL64aeGqbtg6c/x7yS7
ubB8Kw9nBiqcek0onZ1eenfFTR3nnfKceN+B523MSDSWuf68qQ74dMKestcf5wDkQsnG5IIWkk/b
cuAT/jEmxuVoNQi6C3imTDITQbTZxxuWE7kuNWdOKKIWWaDCxma0JZY0tY/onQ3f7ONxFjhjoSwm
+HXq5GE3GVyBfOhLUlHJt21uspoB/rsXhN24uwpn7H5sbsSXrGo/lMJ3pJzAfJoVatfF5irtvLfA
3vpM3InTo106JRYnNsaFI8JUUf6+QRKzIR/9MIr1DPGF+6d2WTcgmzrtH0YjH82wcRmh9QnnTMxy
zVmJOVrfADLbUfygsi6Pfr11q3q/sBLzFu8WcHTfhio9gtIL/2rQq1v2tiA4Mi9IYQ5n0Z09o3gq
pOIV2iH4tVjzauuLBJEQBLq+wgoqbb/1c+HhnQUZ9vfn8bzb4p4vam9CtONHVfBlGXl+JBCuv4q2
xHuRL37ppfXGex5TlGT4xZXUR+tco0jogtqMh+e5VWovqyfyEUKSragx29mtLBycH8qzW6Pxe+5R
XMq08zXKRIyfIIcERwRgZG0oOYxQSvgRf/c1tjCm0vDQajNLLV7XKTQPdCbLDCynT57XpBCJbGLG
Sx3QOUAay8BgjSuOKPvMe3cHjiNMtcu20D8RP7c/EWvYzTJvvPkNW5Jud85YebIWmTbWPDPXhOYt
7zO7OfKcM6E2k91pLl5bKz6kPQi3cLOUKiinSVhbqhPjkr+5XUegH2tf4uebR0PG+HLpt9f45Qvp
xCMsanWyQFSjna60rHrQgqIeBjbepaf2g77+NYZWy3/a4l0gPx2lv9x5edLJacL/M0PUMxDi1+/N
OF+8heRLxyXdoZocE0xc194xobPTqG46Msg9dx6dwg6lIPlKM4zh/yLGA6wT6ICjDA3tJtaP24E8
iP0xsrdjqm5hxcz0B9oZKkOUQ40HTA8q4t4Ie54B1XC8mWTsX8LvjfOhUWtvBNH3rGCzoU/BaLiO
IEtP5zxQK3WSJqfHWMeyE9s9xFH6YqSAxIejSkrEBhmeF9Jv+OF62iBJ2INIbTJnxyTXb7M4r6UP
QMKtp26rl5J32P05KPaFbcyFS5WX+pIkCRuYExDQTbqdFSihpSj9Bao+nq9gA2qRg5KWLeiS/pvJ
v/5kEjjVIo1MGoo5e4GThptUjFCd4G+hJUkl3Tj92vhL9M7epS334SRgh4msHx73YY7emunBqb5K
D7LJTuSlgK2z2bT3D9S5G9tZmAV+2yCS+t0KABX2bKIaJ2KQxy3n09nkLSIUnRUAx7zgWVXwJnRh
M95UrS56wHmHHDSRpxllU/j3Br/kQYyDXZnIeizkNCBXj+C6RCPCSurEUKXqziV8yE7YGTTs2Huu
lcjyvuI8zn1mmw1LVeRn1iotNfMIvuCQS6zj8EP9m7ZJ4qRPfo2cjB6qYX5dTXttC3y/OgHftS+D
cNsA+v6He3dpPnrNnKdJpMeiHbf/IzNs5l77QYoY+cZJT+rZ7RlTyBo0R/CviOOkIn71uatqNesg
BfQkur+4Pddo9lWxp8/J5O7E9Jhy0e3Q+QlIRrGKGcyqyD3hUXtOYkWON1btcSxKM3FELX6+8wBL
RT/T8oUOvxG/eGc+vN79IaoapohYGEzyRRXr5UM1S032u8fndp+86Ba+RFpNM0amfgy1FGup9iBU
ak1fZjgI4+S/pRpRWaZWmI/a5s61z7DlWObohQJSIUyXv/kJ1JXf6SwGhHFaksnDDkLQwEzg9pOu
hk7+aIJvyt3NFwgBxF/ZbiDlmq3ICxm68mbEP9m8tVkYV4r2IWXUAn2MMNtr7TgjJGTWmjF++VjV
ZqR5vVsOUQjKqjycX4PoA56eIuqCLoGVMeT9vOAJ9ZbLrgSWJSOK1eZiYl4tsmHIeIlZZYZWiOnD
Ow8KJhq8E83XStGml8sDfDzx/3/BlO9pOUOAYY99gZc3svVjO58j+9PfjJwv60sqGE+EXufGAynh
xIoFJ6CSar+K1yDy5lWe9DOl5b+UulrDkr0QWZsDSQKY7sQ5lJPowOkZA8LYUZD/63Aq8lbfN4iN
upM2QNIuu3AblJuVwI0KDivqXXRTvgdfyttolcOrD7fMNv6nOqIZY2MPZfcRGa22Pw14p8sIwW7C
wH5pugpScr3A+TleereIInPYFvcS3r3v7wTRlVJvpQTtMQoUY3JjCySEDIhiF9upvrYwOjmno1uo
LifxLZWwlJp/wX1AKS+DH3a9lojl+c4z+UYtk+79EyiPonnOFm2G5yimmxr1O0vMTwuUDE7u2h6/
3irJurZR0gov6QRJF6LwNpLa2WyfCevxJqvg1CeZ6seF61GWeWxI2lLbuTpsOgwgN+qk5O+EoTMn
BWMnN8B+7AtTWhL+00z1oQ5oY2Nl0lXFnYokkj1Rp6k0rHQAhGclEC5jyq2i2xlaa/5Z1DW9BlsV
+GpOatvrY745qDVEtBfQJiLl2pFJqp1IwOwdoL1Qzpf4H8Aef0zDmBqHnKu2hsY8zcmo7Q4YYFeb
+/uwtrqzTrYZ/1spYquHbai93hPPLbNjahzFD8SkZfpB4buG9A1qNuSxsUO2D8X+zjqpKufkPPwk
XrK44wTWXfgaxpeAVCaIEMzkZGkFIgQ2oN4Rnx8lOer2zpcBslKp4QG/xhSg4Q7R7618hv8AhGHb
+5vvQBNReUhzRuBGdIlxHywguLLIadkU3Vj5N9FrYj97RXiPdPHY1XJ4z34uBwjHBhT+52KVLqaP
Q7Rc5qjCl7+1o65gOUQJdCv2KU/6YdEnsXZXpmLfyT96LGmpUROa3HDElNwDfF+yejjBdvm6Ft0R
om+LiIzq5ry/+LUui1FXcxG11MLBVSNJ6BLcGu/sTWdds3OALqJmk+7UD4B4AjqW3v/wIFM0D+tm
dzkOwSp25wH5aXijRu5KkY2BeJpMp/blEwYoE7cppBBPpOnWnuFeG2NNKfI40ROyq/KgenKL8pHd
PHvBcFahDBaZ9yT/ID4/3ielcLGrPGc1GiltuKqAccy9Xh71baDbfpAvks8O2odYpycMcNKuxg+t
rMRcU5D3aC7mgrf6gGxBMc5iOqmULwGcFRK05V0pOPUWprCJONrJkvRkTpo3S/n0eiso+Dcol83Q
Jz3S3IVPpFi1bqn8eOQ8gZuChOIYgi+7FE6mx45j1IlFYF5whrx4NvW7Mb4dAPEtlEEAkKcol55q
DHEOcZSaD6xRHRXkdgVeAIeV2oxcHi8t12/uOdTjHMS/vsPki3oqHKhGu0wt6VUgF7bQH+OLlIKS
qtqWmmz3XDQ66e2f8QUTjc5ft3QdJawNYXxZNAIp+qNigms9NNFnKjpLAyNUxZGXv35UHD+3ij/p
9RWFjmzqVrf+EvBUkHTYg48PXMT/e3G2kLucBmYXEkCuYRaPuOLLsohLMboEROsWoFniYfl13r2g
evdNpmxvzhWSSdzFLMKvwYyWM8GfD72RTfR8Z+Nf8i0oKbjJ0sQl+n8rPTDiEoeCBt9vg0DKzr9m
PCmLVZN/OuYq5jxQfAkmmVlNh0PcHeYaCASYhN5vgh1lxJBrUPinq6rgPEuYPZRXK2PVrIaIOki1
dOU9PY7Cs8m66rMqsMyMmoJP4oSbijvs1s3Bvx8ha/ybctmx1ukN66OFea+CUaJm2NohGxaq8E97
dX0cp6muYgiT6rcGZ04M5OZs+zDcCD3NDOHaB+lewz7VNGUwQGnaWwU65QPORNRaBAqNm20L9RQ1
iYp3sLNBz7yG3iNIuZDfMolaIfuILFE2P7aYCWerK9Lhv8n0JiY+x4cRo9ICa+WCnqlvZu0OUmOT
KMv73gV8vEjeiRwatLLSBHNuitSOkAEhM1ZWZi6z8yn779csH/N8HoX3VCLWZhmiZxfdaM27Yeuo
dPcntJF7EUyfaz86+2UvLvOPJTh9DWu04ahZuPR5oczuhqpRaqRX4wEWPkPKXXwX70RthYfGbU7G
kKyZk+WQLj25iiEbUHxKu7uAdrBXIAys90+kHrA8AZHfmKslzQdBMY0+oVikHlxcQ80uS4hKRvaJ
KhL7gdm3OgrcxMzwcSpq7C920Ul1S7XTa36olvIg+XQgSvs58dsn/ZzRHTE1xsUTq7W7EtMIIk35
unGoJUf/fgqb34i2kyh8L5GeY0c6HewCtDdzCMbdlIRx4FfD1J13Qdi+2ej2elgcr1FfDwKeusRC
fPPg8rlmGXkxoJUSOkI2f9ukBAKJ19N5Z2WjVD1DKeIn1ztDKjz8emglZzI3/SvQOddThgaNVEhV
k9Z8EF/aFR0Abu0tbDQrAap+gpdDA9aULN/939PCkgkL1BV/W3rYGrfz+NAEJOTqBUHx3RuXJgWl
LwmAHuwx8VlN7q7wag+mDyfc+xJ4ajHgDTS4RvF5HRgBgG0+2Pnejy5PIX9W2mdzLC9v0lq6kvxP
JRvNJRaG8pAGyUd6Tl6A4Y3KXRWw7HCCAzAtib2OvjyGnf2KO0ag8UGfD2/K3FHP/0SqMX2ijVbo
16n8TflUu0pzSLUZ3gFipi8hpzsi0JK1tadsKK9Lp8vCuhIlOMcl0Hw+I4RkMTIuJbjUhY1NZ/gG
WSgLP0dGeoGZvBZIIlZmi/MxECvNS1y1f0jKCNQ5O5FK98NJw78/50ijIVUfXSM8RWG8vneajFO9
+CTVCFKjzAvF3p0M3DCePwmv7ySqjD/bg5aCqNzLclDybFLUdF2vrqjrqqsr3jK3M06FwOrOU7Gv
ZKyL1PzSm74bhSaNpe+9EtAO2ncet1MhnNwhlq0fx0Xh0EiznAQVU2gUgdztUPXbs4EkqikeQuik
sUwMDbrvXXkJtAoBX06cIAXuP3oSJ9BQsN0FGtVL9OikaYW96DCxyO6prjz7KFnBoXkuWnnhcaqo
fi9cT6vcFp1ImT/2V+OtFAnllQk+xB+KXhcPrSRlb7TbRxi5WM+sn/xkCicvsD5KKMnWlzuQHzzX
ZKVUiE+AwQsZVRShRxMpn/VOizMGf0prEGgrgug5DddMR926+dky8dcL7ru/fCVD3dLXhJbfL8Wl
1gt5H1ZCmgQzXKdAuMLxn6NgdtGZ3V7JaQJ3KRxgXkFNFbNtio85IDBueJLEH3ANnRXwqV1H68ph
sg/69bzVP3kJbKAS3++ijgNXJvz3TayKfi5g/3+47HH155Pf/MtN+cejiyn2criwdqjzHstlBB8F
xbK9Cg/wFGWUw8ELtj3PSUfWEBfjkv+HeOGES9JrP6o6pEPjOkeF30dUKmB/O7FwGntpwN6RWdTB
rYHsg/OgU01Uqb/ibmEdudh/lbl0Y/rhXXZSGYh9o4ni2A0+NrF6VGA3mXcuhUyHxX96Ldg+8MVr
tjGZT6WqTV3sH2fbksyhCFzTfhnnNQrBzg28QBOtj3+9HdMFlzJzvKb9j/LWNUSFD10Wh51GsHB2
ocMfX7eaf7BSrHfia0Ee01tAJIMxpCxZeYPGYkyzXF1dEITTD3r7DD1Y/Pz+qz7+kTlEYD/s2GCW
kiUEOdkX1pDmutCrPLxo6LxmMyqEh3oIpEH1E6+YmOBhy1bnxJGK2gSuTLgeKVIuuV02wApH2JHM
nGL5FI/wEea0uoYKPJ9yuWNy/a8aqum8k2a6EUAniMfiYCicQa3DzU82HuF/IIvwgH2u19CGyAgt
aBVM4qvA7JCFB3xSd0G2Kolejl1hcus9XYF07sg0uywlsnObycZ5KQ7K9oFZ36S12T2QNrOTv9Cd
9tKDQ9ZSJd+yMPhrRLV0ZTAgJKEzH2OuC/6GGHtWPpiLi3nX7OB5CTffJottbWAZdId2dWWPBvcB
tJOY5uoAp/6K4b1NnW4iapUZ24O9wc7UXvJI4tAq/7hlUNbV5TMwST0trchgrxhzFstdCB8Lahsx
eT4I2JaAXH0Vo7ssAo/Dk5itWhRhktRHhME4gSuhR0mfPjCykwlojzdOlatAm/U4kHkkeqSOKMmQ
9PSRt6TJOOVCE33X4acZ0XAVygnq7Gc0bGG3d8rbm+Iklplh0nyesSn4LXq5+HXgwNPsBCFDd0Tv
e55AciF6fhK3eZbVeuBj0dVyTKKTGUYMP4blZZE+V3apU3O2fuCac4NCQAeHPL24AanoWGBzO5aA
KCoTKVysBlvzlhdcDSvBvoI4QU4LNDVAndq0KN10/3Q+l4l9WK5siZr8xGfUORJutVTUyZZfy9LL
Cx+6gGA/ra9SvIR8Jo8vaaZvKG2kjO29D3ntoJtglWYSsEOCiy+TIw2sSMcL/HjEa3Z5G05N3SgG
LqGOfO7UQh6dkGuOFriDBUnIOztqfLN8NlwlGWCFoQ82uJb5A5NUNPd6Yx9e/pN+PTmw7vS9tYm1
qV0M143TrujgB2W5wjv/6JL1G90F0rkfVQFRXNjJklxObdUK7APIDuDn7KQMQQJ27gMSRF/vpUDx
ilWtlb6v65wBwFUoPEKT3Q4DYSW7VkwvIEaeB2KLZH+W3WnUk37TThtyXeJkZ8EIdxq7Kj9R3x6u
p3jwuBZPLdLINPtuufJbXQFhOzawHL5XhyseBoDYCH2OdqEWf7WGLPKdQuEzUAARcmqn3R28LmUk
8e9o3+lcMMohqeh6xKIZTBqLzvw9NvQUjdF2/YLipFdkdNh+skxlR6hkKJtf6oIUED5+0erTxKzo
Z+/SsyMER9zXZcbvMbFLnGQ8D7CzcgK+WKvAttGZ9ckN9A9dZDgXHTHscMc5B1rDQcdHOpploFZ1
vbnClnn7GT6bbSZKpvOSoFymlFv1DQOo8sE1JHxnlZ9WhKxZY9cxtpy1GN2nCrRhZ+M3cT8OTGBZ
1kX7XdArffDxNkbxiT1gm8t7KfShipRKgUGlUS8ZF4j+ICV4LYgwNjpS+lpMUxRN1eLxQQ3Dq3s7
3ALEbg54ssanBfGw9paRinkJL+BqkAiZa89rxaZMF0M8Hg8Lmm7v8LKchvVQAaeLhN/y3SLYDZ6W
1oWMtlyckbcSPdT6emEKJAeYVm2LxemMG9WHBaIIJhyVOGs2C6KWE+GO4UL4Ik20c4fDxzd8VeGi
ePdQFctEhUTGjrspsGk2tqxGpJHoWTEFcBCv/43/2JLlOGB7YtEdDlpONFvvgVjfks8m5k5sE876
GVV/LAMgb6OQSSlL9m7hAHDhR+yc7Q90nWQDUuSkj8W0bGWaJU//q5TftfOQu1y/XpTAXpLnjEZ5
xjOouSgSu9H+f3vkxnOFMLP+lAnqt/L0jSWUdVyMGFH6rgjH+hslbkHg24IcBoRK05YGxWg5drea
tu+wBH7IWfaPsxV8X2XPp/5NCIciyXgxh8b1SHcsgSFky3kB9GKW4o9CN58thm6boChMVlai+7tL
LNgJs6ScQnGKWrMb3+OJ9bvm+4ge3dkK7NDJOodQ3vVAMm/noB6EWPqAwAa5VfmsngLk+UvW5hPl
po1Ku6qcPkMPy8e9kmmwpVSM6PgQwrHGv98VyqZ1mgbBAL3Cv4itWWdTqHwXhJFMwtYN4DAEROY/
JsBRCOOWepGLS5oj4n0AQ6tGXMluTsCQ1iEud6pwdrH0UKNnU2fDfkP8VcYLwuir9lePTIVaqear
wR/1OownyuyTAy6r9tYw3dI3kdmNPxAgmcJAmtKdmwhapIJsqR1H3PKs5KVCwoK5PzRQhMgEcjx0
8aUvDCarn4ytkWNzZT176a2EsP4fZVPF7I7nNhkF6WQ3mnX4fGZBrcwq6GPJq2mQm+eiQnNtYDqO
4tksXP7G0lTN1DyEU+cjDWWjrvYSiUeIVkQ8tcg9CJMqMoXl1ovyQpJYJiLV4xsLiLfvMeGdlHEM
hi+lylpAWedaEt75Y5HmkFSjZQyyFYi+iFcKLgKeyTYpoM6/KNMLJo5H5mjOj094Mo6pQFrYvhSL
jSKyG6kP86q0tevu7LBiQdZzUrZvvOAXnvC3Df8KaCR6WvFIZp134piOC9fnXuhVBHGUiZ8tWRiX
QNCtVdZEpOisVdde/IsFA2lXah89t281Va6Iwf+vMCZE6lz2ns5R8ZLrEVL8hB/86n64U1orxTAU
bBYnlXZEc45G/A1vvHlt7xqzDfsqyoVxBbS01ZS0S2DQjcA5HIfRVsgOy6JOxLGuJpKmZbXgMhWo
3zc/Uk7Ol/Ce3nhZBKQx9048aaskMySumPPLXXQMKo9mVuqof7sImuwyHtHkeidY86Hc8IQfpi/W
/wF3l73nXpOBf3K6e6sAl+wxf1nVrNPrP5GXAQfD2kjedf4FFrMjM7pBy+R4Lo421rADFyDDSJ6Q
1oI6BB0IL0v9L5xaNgl+2lG9O8hFh0Ir3O2bbYjI7Tu8MSW7A0/xBWcXkNGn1RJ0yD9K/4xZiErR
Z9Qaaiz2FUOiVXbsGEBjT0FzR7sXD4aPraU5y/zwyzcGGNrsfPmZYECQhVDNK3Wz1fULf9KaDUNo
+ETLddknk9Vfl/iKKDVdd8MAVBiKZnxxztYvDh8Qz1IvUHzZbMROyGbpcXhFdKNzBDAXe4oc5eNR
EDEREMgFWomwgmXReHRPj9yeJ+ywroYQG0Fe+RDJJqvDOFkTHipnMC6g8vJVdMcMQvAJK/Xe8N0d
AuAkGYoSFo8s47VXhtHRAzm5xoURfU/jpWzDci1o0Qw4J9vYM+y4H5qQebsCW9uYu/78vhTb6YFI
+vs5XiiJpvGhz0Ooeo13XAm5BFmGmV5EbwUEh9NrTaZRbch20WefLkvT7xKgQPNN7UcpzVHZgAhp
zh0e2hCNiPj0G3vdWwT6fPFqKtMsr8kWM2P3D+utry/3Giftvr6I4DqKRPzf68getQgRn0R+sJ7g
AzPu8K5cQCUHTq13LG7unM7cuuHsMADPqLUOxl55R1EWm9NjNjnq16wUsLMn0ck/NF5fB/+uhgMC
kBlpJONRYxzlkCnClNsXh1kYD1fyDi7cH+zHz5RMj2WRrKui8ayxptZ27tQcX5+oK94STQtl9MXm
EGbhu3UZISIEgUXzsdmhpGWw6+NbQo02yuibVjo+CEqr9oiRSJLiuRcn1BWzQSYbESmKYA/jQ82n
gnNHr1na+kPqkFtFpujgoTOlFGvAP/pb2eOEXD1nsCYxjPw/dgw3wIR6xxEoYUlLxTf2unoLr6Ew
ZMITzKIUcD+BYLksGtwi3KDK6sNPqiHRi1HUQdY5geUhAU42blDc3v+XzFEwMh6/PEzwRmj7RD7i
eJJsEn9/WsNwZ8g5Qu2VwaNaf3nBOzjuPO/ex6L1SJHVo7xI3b0sGxMaE/SA8Md89VBXMWa0Gck5
4wJGzr2k8GFJZG9UeWYwOyCkujHXfE/aEq41qrop6/Uh5exJ1XiEiT/QDx5sSAtRZMNVy/Rwq/qw
EFgTblsCVZd5s2ZixtjXp5+RtAz1tZ5oFPnpjjj5hw0p+9hevt0xHIeGWa6LHGPxplSEcWlNrZeK
fpxvqyhH4FreaX5JmDqGzO8JnmYXxghLGVaPMxQjHXlwOdia8pprepFmp7HzEP8+lZv10AKsrGKz
dGGt9uYJVSVvxUz6dGBk14dMdUDbx0jXxe/g4LaOZ75HYaaHln7ZfHMCEcMf1zvlGNA+UTF+akE1
SdQaEYvQtcnPRGllzyNPqnjEov+H1nFwwS1wi/7w520WJsuOllJzE0ss9W2RtPdb6bcVxjMD7NKF
X8wNyuK2YhvQ7E3bwQSbtJSHizeTkhavZ6Tb/WXMGdVUVQlejxsrtt9tJuvkZwNzKgRK/cFv4iVS
GFOeseFkUdpz/hmWUmBvN4SxhcZhdi+uC7xvfDDjlD0tCh6qcIAEM6TyHumj26omEgeoBbwk9mJe
3uxlMGiszjzBzfRlvXozyQiXujfhcCmQxwC8/3uKaB/nvRyRieM9IMiD867ELgtFiZAQROEAIHmu
y6PuhVH4UBw2OWpmocDrB1e/XFB4eGQDmY2f4YFLNzARiw/zjBDDOL4uflGB/wjh6zfZvi/m4QXx
WKACNsMNlQDNM9Rc5V913Umkc2wgNIgv3+6bbBNzscdoa7U3G4Q/KIPuE119PPgxzj2rE21XA7tz
/PWchyBbvv1S/m3AKgV2UvgmXME1Or8+I0jFHewsh8qOzj1fDQezZ6pCNMGpQAccTqYZW1wjhIFc
HuXgjczXsuLybex9ECOUpEoiyJQXw05LibE+oSE+D0mp6hbGXCQBH2zzh00LR0nWTuOVpMjOMNiZ
+eXtbd6Lf202U/YKaa4I63LitCi94jCqTGGXW3qxCjY8c85zo/M2rIIDk8KWaHY9mYX4FZl59ehU
DaC6kwtVg56QPftGmJTqBcCSYzNE7xFDbOKgoZcuE5T1RFsZ0/ThDXc0vaCuLlHVqBmWUtY7t3OU
QOXcrCQsg75CDnjPv/9Zw+oUIqNQIauSI5fl92uGVIKoEhVkg3RjITjcwd066qeCs3gS5b7lcGx0
rzeWZINXlXltokuloZYz2e34XbOQolvuoZJAUVzR4wgwlrKg9Rqmf6DPpFttbwjvNxT9qoxHibIa
5e2R3y64r5xHySFIU83VDHyRywdEQyBKbHeae3zT9ugdamilPu/67tUMGzlBN1Bi0YBCHcg8lqvD
Zpku81UQU18iI98Cb78qm0MigZrJHMZpy0oiIQcEi6tsIeX51K/j1S+VFAaWQXKTb9OfxO27lvU/
sbcFvAkX8J3Ew1lnVwV/jhkalDdpwGAR0YOfUKTfYE+rG/IGji/7xcx2KhSQm8WMPO42WLEnUTXP
bEA0Ya9bqCDc1thswrY9yfaX51ReaaiE1BJscA7rM43a29nJiEFPabMrOFiJ+7bhJ2aBEybI2NyP
HcoH6bELSr//y2LOlOeUt+kD84HUpOw7ljHLrQqQkKwqfMM9Nc9T/ZaLrxfhngRr/x2+W00hjZve
UdK99sprEdQS/0MJeXj+EB3fLLVcRxj2lZsdsanEExXeFnovBJKs5ATOiRJPoibq4wci0grAHVfh
/WBgcbKqrb13kkA1NKTUQIpmyBS+a50g+wk2AkAxHCyVjf5MTiyaUjVrHSvHNEm6ZhVjKfacy5+N
kA0FvYKnQr+gr8y9UewGLepcBcWtbzAgUzPF822x6Hi6ISWnHMnjSiW7mudJWYiHzqmY0+VAvby4
dNkOZcKwFWDs1EYOBYk5BZTkaaT0gxvviTF0ogUIY7Zb7w2EhTl0WU58iEOQbGint3lmBlkl8mmZ
zz4Kixhjxtz6qzMbHOEEiSE0qVOv0s4evwTrMUXAtKUKCc2kQkPD6OQRL3OlIDm3BZSLkHqONBvj
vvDrBC7/izHf/1YW7ntGdxnIgiHHmzinxuFHrqSVsjOntqaIuywLovQ2s6VJzORZnGAAeAMAkBtw
6BDm/+Bp89XyTZSQMMJ5uN4xYEZAdKwHfrnYZszQMN78IwqaWD6DQ5oMe+e4UsBBR3VqDSL5yzGY
XpnsSmRc6pyzkLnpJdLjN1w+uAWkeBbEUGDip7Arpb7QwR4gaa0vaFqtHWWvP7ft1dWlz3uhag0K
k6doIF4iD4xPmGQFGEEoBXfhPbjyTJn4ZwJyrBOQa8Gv07f1UjeUHpWFPU44HDEb1vuzeZfhePgp
YuLIDxduxm3N+FK2pvpcNx1ge0CmT3iX5Up30NKipcnhMxPSSQ7UZSaem8mBOxBRK0naGK68nJnn
0Roo7eapVnuN7wp7CZ51hxE3oD3jtXC7AeebkwmlHDtVtGF6EMS6cIPTCnh3CWWmLOL/EHnmi790
OmxeR/3wFNsoGP12Wwp37I5dOm4ORv76nltk4zxCR7qNmUvAYvNLPyWdffD9JZnGbjSCZEyK2tXl
wxoPPEEbyTUpesim1WScDIDSeSnc7PEg6hWwKFitAh86+owOjyOvWxvS8nk0QmRi9blawJhn1yoa
EQK0YyHCnWcjggXwFtTVSZfyvD+YTLCQ/hXQMq2T7yXKBfazp9O9Xtu/m6Q2mLDaFG+CjIJb15j8
p458KwwnWiLQy+IFYqzNf/ihd97+2UV1rQuw0D+lUSD4+ALQd4RWcRMVqAdu0xi2d0Foa5l28Vk5
n2zxsNWEgYS5oES6jW2w1S7YuPZ82QBQSlP2Mi2QJUxzl/B4p+B28wP5w4bbQ5AtCbIJLCgOKMua
s1qlecfc+X4IVOtyxfFFU/q7uPSrp88kZtrvkkR26BsJNymkJqFXTOU6J3HU1pnXKJGPLFKvQkTB
4+4WLxKlA1rZOtFl8G1QnSmG3UJ5OAtIHRUuvgrSuVqfHc/oRQ1E+K4aYVzObWhGSOuaxM5wj+nV
Fa7u5QHYfAjTdnGxou5grPcFxx//HN4mJGqo7rrw4iEWm7wIsBtavhLJCyvBh0r7QHcd4CSjX8dm
d1kGolIKlZZbQwKRghvTL3/ylMd5Aj6SFd4LAYB2OnIC3r4hJvtSM29zTX5kC2MdCbbggyGqhigB
8JqAaZgO660BpEOhO0+um0sHmoSHT77I1MxGV4ma4sB2s4uN8/Y6oTUAYMIza6qTvXqM7MxalGC/
MOTGqV8Cyx0rq6a5QjiaQgIrd9lkZ5aBGXyFxyDd7mjFlw0w7VKUmgNAwm0+9CLMxhjoPhHQnpNC
jK84UBtFCTmDnpRMgiR3cXUqYZDtVi168JJnCxeJniTlEp7pfnylypGzfWvXR3jX8nPvtU4MWM3+
LSCpfVT0JJmTMeRdUd/VCrSuV+RARzEYv9XtJsfFS0Hah/b8FUZH2QMUT0VQAkmMJvKl2agusRsR
O0rKVq32JB2mbjCcGJdnX1mrUTMwX6lyoyzC1qOgXynGcogzwjeuoqaOl+ZbZf2kXLpp7jveXs7R
qYrDG9TuAt/asMiautPmiLgqfi1fB8hycqQgA4qdUpdJMjeTbJPUA3r8wADYG3tLQ7VLYMqAe/qA
nwlYb0JvK6Uz+/FXYbRCNaqDi6q5idHynRfVWTulkvlEf66qBwMoZ5peL1oEbbJ63aQX7wXNVkjX
sZOfMx2jk17sFeAwZQUpiF0ORKJu0hs0c+dnmfV2gxTmBiIzOIMZGR+3HZS4PaF5wGQWo+EV66KK
k6YyFQGBEP7FBV2zRW0nzLvTQGeVoiPytouiWcAfj3dywbg6aB44uWn/QMobq82HrZ5jPu/+0fFA
+0euErrjn0CjFue8u0/6O16Z1qozAkiERN+RaKzY9xrfslH9PiAzvrLgxRoNw+g0HN570qfuNUMB
w41Urwz4AErb3u4D2OV8+uZHTnyite775ZJTFmYpUs5eOOmMUfL1PunumX3eEMcZPrJUco9bOFuj
AXYJc3FCSuhJEoHWWrYcIMBKUWjkZENyNfJxbww22b5Hp5GAnkb/yvzqIiTi2wHID0pDZQ6qTW4m
fBxdDxpf5xU9/V+4iqEtgbRlNRw4NmHVCGAKH3HN2w/K1Qn0NoELVPBK1mXYWwBQOPEQK6o1TJ+C
V5KgaMyJDAYMxRUfCVk03LX1edRkUY/OLOLHQ7yItDY9p9/ETGrI6wvk8gIJGQ1KGyWikbZIvYW8
DcnlPEMn37jJYNP09s2FFeaf5GgEVUaWkavUC4ZNf1BsSMLU8hzAZOppWZS8iDASBkzfQSWvOmm5
/EcY/TyN/QPzk30WBXXuPhreeRIN05aRhU6U5Vm+P7rIdV7C4/pDpCpiM0SpJeTtTgsTECG8D/8u
XWsnEwumpCbjTvHZnDEoRGjbIgmJgqNNLzK9PzQBFO0yhwcjvGj/NRIhK90SODkroDTzp+qB4kwu
baS9fwEQ4ABhKKwrSn8dfXhEaSrsXrofwhImAW5Gz/Gx2Wc+DZrY3v46P8TWuKab0bwVLWv65GQC
MxjrpZrvqEBqUHxbiV+o+nvbHnHWXUehHN1VPm5C3ptuil/fkl4yWd+XWD9TL2H/ZmH/BVq2HuMx
6hmf8IFAnXpEq4Fe6rkbASPM4t1JlOvNaXgm1JByzYTf5yyeExjR/GtahB24SVvjNYhQ01/BVo+C
7H2QWL2YM+/RvMUYJNNVfOWWOKAm82PaQDs4ccC+FO7uN8agjVhz2ZRJ85P6LLn4+zgatmnNxYhp
EsBuICbvaM7JQ+crEQuANA0ypzDGSOPxQWdPG0EVh1likzZB1kFfqqcHaW4d9H+8xDDxv+PP0lFY
1iKql7eXSHrBrgkz2QBC10ATTGG2gnp89nqwO3BRGn7c0e+b+zheRniAvJjsA8fdJpUzgF4vGVnn
1HoNUyopNBd0YfhaAoE8D2HHGq6S9bvuvPQtG+kCA5h8VXMWlWCw/WOpRgqBdmh6S3VVu5uz8/yT
JTnSkn1ehBAhr0uUYr7Yj9w0yjzZnpjMUC2J43odN/44bW4yze4KVb4V3OU8gnqklAabyL6BKScs
kcwfjD7FgeXaME/b2AGqCuRObyvOaIXUlXxYyhVttzkopcaN2sZB3ZGFrv51fkpgF0Oedzpswe7b
mqFRiQIDTY0NvdxcRj4ULjFAz+dp2rIBj6thpD6//vrqzgMk6Rv2AoBiI9kQ4znkGqwk3A+exJIx
lB+KUl56jqJmqd+11voaS9j/9fFnyI4ggeVqeor7QCqRWA35ja0drlSUVv4E3bE+IU/UnaRrUI1s
T8fc6j3qLhREvsz28cy/l7gwvtU+roOB1wzDxg4z6z+AYTWNbgASctfkWMcsdSB6p1KVGTF1gopt
dc64GVRut9omLkpJPm3FU3jab/jAVE77TSvGUsTMK1ZBimqPYNZ1oLaRldVNllq0hxXezAygnO0P
feNEG3f+KOOqv7vT10AYFdo6uEbMvYCyE/afc1/n9h1xr339IA/weecJ9F0xX31pO9N70YjElCRC
lXDRrM/yDghUOeL/hqLP0iX0U3UuWb80OJiIKAgjJ40UjyQOYoQxLTUW1BmL1sfnYerefhk2YuYc
CW71sBBqiIlyjXNGMC+RX9y6ErNw3V6218A7SeOZ5uTfOHdHz9nVCwXC1bdK/cJWGQDJVqE09OMC
Rx/hDICtn6G1je1i35wEtdZ3hb3toebN7rrOv+c2UVvQBIqzqifYZofXU+ucRP67KvvXTwCLzfa9
ED33HiDroLDRXndZdYR35Y7nifFLuN+2Q6upP+UEYrMVHGvSes08aihkJO4PewYIll63iZDM5NiQ
VPLDu6dt/XQ3+k4YFCY7UyJD0tY1bVzf+eRRsx+lvUodb/n2eGkwmRMSeFPZV2VGh3hLSWw8MGQk
NsHmniaky0sBGLiv+mXxWp/gcuqs0rEqgL6lNJjI5Ap9hNNCrZUBGJvHhBcPWmu7ChDfG+ogjenN
5HQYTqtjVRuvZ0/sVWhYddwxMJOQHaToUcmlzKMaqZjToYc+XjfMmyzn8zxGTBgrrzpApijxjgON
+xpj8EYqVAOo9qEyBXZUkX5zMAIn+/OGv8Z3U9RYRsJOeLuhdnT1bXQ0bq6B8OVMt4mwyezD32i3
luOpscMeR+hRtDwraHcmiPuzO2HXb6ymNdvIgkSZBZ9cKuQpCGd9w+pLSmxkesKBaV4hnbx7sAfW
a0SL0lpS2jNLyd63DBzJplKugxLw4RbKWT143OYRFJ4znNEzpoulbXhV9vh0wQk4axYLupAR3z0b
ihlsVNqMlEQxN7bAoeFaiSmBrqC68LK0K11DwJucMWL0fLOZefUSXNwwsT5SS2mwGD0mbdkuhjCx
/SmigWT1+qsaG+v6VjzEEPgSFPHR22uG/ubGPx115b1XoxPRYMq3KR/F7FyErwiI/g4jvv4bh/6o
ueUTksHTN71SZHA5+TLLTAjsGVs8OO8GT2qnRL5UyV0X/YLq7ZbPdZYH3oCbiKpvBLvC71bxSw8H
mjI4IYrRTlqRdc4O+MqFyaobysjrDsHkGp/VgZBDWOx3jjnwb0ftZzQva7Fr6ls3M52pf2aVvNLG
Sk7WZFppv0rqyus+lNJd15G8YV22qdmri6plJZSBeqpckoAuXG5JgrksFKeBRnKJdsL5OUqJSBve
xyHPDW9olZUfSW6Igpo+a1d7mWey9ZphmiAIj48xKpWcqdWU7iV8VQs2ihrIPwOsuLbUNr4jLf6t
QPzclywE+iTLEoI9de8I7gY1B8p1eoFDvUmMfYPrx5caTkNWeT/4J01u+jIHSOXoKpWGxQ+xpqgD
2E0CUjsacnKGlIw66d8JZMG7/nwzrt7TC4QLtKJPCi05R0B4GKQV99bzzmAcI0nRUh30y4RNErsk
WN8IP+5tkvRWyeNjUkneiqGUsYKbHdvMLklNA1VzixdFFgBXo8P6ziT5h5P7w8jK+jGrtcmWhJxn
3SAwGEdPKpAuVkwvLKd804WHdg+Nn5CE0fJUXNGVEu5FqnwkAqDwrplwwW/DwhZ9WQzx6WOSmVK+
yNNnrUn13181+J3LCgQVxxEw36NMQfmoPyeZUQtzTzO0+8P/X0q4YWOnsjh1L4+sUI8FnC3VHv+7
gDq0TRsuLZt7rfzA3rqiEltPUf5+J3CJ6gAD5Z9z6MPIRKiIYSs2nDdMP10/NkN+qyxxEIItnLB6
j7uiOyOemc2A4dsNZhrzUvHq6IJFkJsO+4FRr0iOpFfMD6uPWF02ripkFNKA0ef+TurDLot6obj6
GVENm4S8HaZljsJ4tSjHZPfW5ALIhemKaCrxLZ6m5cPveMCgfrBFsBNYy7JHgqDcCInC1W0R5RSk
7Dw/Cl/rCjNDROf8iHSFwya3eiAs7Pij1mjBAlPg5T/hau5P14HSQkC41fZHneqmA5M5EqfrIzOY
Oe5PQog4gPPPHsG7Gw8whw1gX/LNjPrlv9aEB2iNCtzPngRr3ZDbE0TWKSM/hIDnxMNwhxxXfsVe
gMc764N3Fkeg7Q8GdIEgyYiOPc9GRUCE1TSToR6cERimP87fIOJ0dlv0Y/nVTS9zc8NcG1qKgtPb
e0oqD3z66QBN4ogte/F/1RliJDGkrPCL+h7uS+Eym16iaDTECsPGainMN7PjXzQATArfXsMh6uHU
hVFxSlGUJBbv/R8FIddrPdUZ2S7LklXVDYpxSz3x9v86BtLGWnoff7q1WJ+2/sQeVecrCOsXIRSu
tGf8OhsORUOAwkiofQY6OpIKZAA5KuFKTyO9lWq8VUXJXAiDg+y2cEi/GwiESQWR5glLdi0YvOmo
t0p8F+srlLTAo/QGrXkBPvggfsbJWSoK1ya76ob3s+tHhPSlBDRcInZTAT57WHgo6nDWjSR3n7fY
NC5hg+i10oFexMbD3cnm2d/g1fO8WuJru+BKeRsf/wJrE1NT94JuM0+d8Advpvd80e42BVziqeGQ
O0ZL9Ww1EJQcsguLP7Bkb8QUWFLkLz5O2W2WX94lyArCCxPBU9lJmW0tIS84KO5akrQ6N4mHP59G
SAO15QmYGMaIjUfPj9Ul0MGaOnGnMr7SAk/+J2//LXUFNH1ytpYIrxLEfZjaR203Oz1y2gzVV4Pd
Py5dVu9F3NjcwP5PJvkptMoFAQiDUq0XzYIfavOJ3bFYqKdFnEHUGbKIHJYafFIzTdk5UAZgamxj
RgtcDqJCGixP5H6XEOoIa1nLqffUG72Y9XGyJ7ajQCW37q6VxLvL/noJLQZVEyrkzehZdx9ITd/w
V20nFqG6DcWRCF+ZpA2NKME7U2lXlB1EHCLPjnLv8GAf7RDcF55XE+Hv/imKa8sBNzFrFazyfJtZ
TLBFuRkVr8K1TGLEkejJPtuIQb/d6TasVlpHk1zJfz3wUWY+F6SOXTrLQ0bFq5Y4JyZz57h3Spa8
FN8kMbr/8e62iRg41Xa2k8o7OgLnVSQFnRn0aUQvxsGsaWzchA8dixsahjxfzHc7mZhoupVAy2kC
KvN6TJtvdcLjgkhOy71iO4oK/qHRXKETSMzdsonwjtNcx/Oq5jQgjOXvlnDrPXkPf+E6qEkTIest
haAf9h/wJ9VIWUolFEdmyJWLAlPXkhoNwn2jmWcQxD22bX+pJTaOjcpEryJ6qHnsX8fopDwyxesl
8Di4PGWXrsqWbZWrGlsuzAyFt1VDU+IVgptjf1L5fIGI/dP9yFY3+Rwc7RUgmjGwavJlRLGjrPsV
2IoQODG9sXg3xGv/aDhJukcxH/PKsZsyP8lvQsLVaAWIfVZTeBhMnCdyImQn2Rd9gRy+n9lG5r5H
cbGxkRlWz8gSarXddXQ/xrOOtw4dLwSLHqQOF8TBBR9JJnVAFnu2xv58TVRKa79tbYatlOGBEwC1
qdKip9Zl2BWkDnWxJYOts+JXZ2Rp1rgAe1NDNzeji+IoTJzkZfp9s0GVPY/5RI0OssBK/sXwCPQ3
8KdLPT1pTxp+xeQZ66XEDkekPl8JeSiJXe+U1+Tllzyy7v49ZlVlSypfYEku04o5/bZVD/m8k+ak
vmeZ1nYynMeOnbFPVw/OH/3aJS95B84/QD6HUu/1pCkq9CIgf1vwtSp6Y9f/uwtZIBKPXT5Crg9h
tRwF4y/D3tKJSswT8pHLVo6HsF/u1oxp9NPLmoNu5vmnAJ/D1LNUrYHcSs8ev31dsbwISKZDDBch
efTuPNuvF2MssCVaJbSFUdDnhSphzLan88sTgGVbG2zP8xZbWuM0DTo7/ahTYOcVyj7Wn5m8McgS
YDF9WFZKXtcfsOj8OpkIYkqSqQ3DNElTAG8ByJgWXhyN7rtSHfS/sqy1cBFlLKyiMm8fQhcF1XYh
Bz4U7aKpkcQjSc53WYdpHZsj+PxTCLrDNvNVwsLjsEVBvWl0MkVTTrVZGUPqhKlGbEm/CE5WXZeQ
Tlaa/bDdZBjs2bdzFxcToiQoOnJe4H2fAqny5ezFgNK1iBFg8fZ/igClInkCl4IS6rbHBeJDH2qk
JhD1KanvXXvJ3LfsE/NLDDdU2KNjyHi81i7iWverjLJIBhC9IR3IZhaLJM9DgoimZR00DrL9c3+U
M3WYtlLFiJZuMZ+J2WNcf8BYEnq6jPA4L/eE8XdclM4TI8KJBQElM2KXhastov+0uZy35+3UYiHh
Zx9wwyJKEtAl02hMjDBKTDUsEWz6LMk43Y0HcfmJvMvZ5mfo0AqtXxBYIstieojBw1PMDbtQx6jD
RGtP6xr+RXGTTxl7hIAoL33dHXCsth74KG3UVzhrqUDq69jTQpc4N6pkF3Map/HBcilAgbmCGa8e
hVokys8/+pyw9d/bxZwT6yOQtZsYQs3Y8r5qB3yCdsOl8UUBCelfcmFQrct/bzyCh/tfP8IrJqgO
FBAnC8ZZy2AcjIvkCGzX62IIlZhroHRXZP6XoIq5iJAp2eLc/Y1+PFfNuaixA4+PGXdzzzTo6OGv
HzcHfAi5NU3ZoZmc5OKTOKfe3ml2OBuOFBGov5loJfay9ly20EAgqm8qiigKN+raXB24h4BAWAJx
FNcrFH2mxYL1er43EZznvI/sb9lcz6adqlJmgdiLmIWfcoGtuHjcl/qy2Cy1+sX/k+QVl3g3m3Ce
AMqVVstgVWbo/bAZvbbE7wXc9TfpCgLUDOlXf4uKQdvcNYiyoXFKl1mRjJ0mvagveBVEGL9Y4sTU
SRyR0C9+L4GXBTyUe53AeZuqLMJdx0miIIHuIqS/Ui358K1v8RGi9apl0ub8SkKFMrpTJJUUh2uN
tlQ1ZrfxO42Xv9JdFHBRPtl6nbZq/WeT4KqwVhVER8DWHAE7J94MKrWkaQVodg4EhGR3QEbpF6Kv
eV8PPSTMjLqg41zDL8bcqeWGQdu46e35o+wXwrqGS3ZrhbTxn/C64lAlSvAX8DY/x5hE8DJPiTKI
07ImOmVMTsBEGBEfKJB1XKUQhToqHohEmXz4Jk4qCkLQ7OFTA/aFrJazg5mz41goyg3wOK1AuOYD
S53FNH7cFGsXwd9f3P7Nognd/Qxnrs7DoyltmkU6axKSN139ZitaQ5WT79FDhvmpSDR0VpFE6n5s
PdQC0T+X7/7x8vR35N5Tf2NblTOgQOHwB/rV+JiAHBR02D5iV4vYZiAu0TAbun6DiPV0xDCTTDkH
lbwZ1EoiL0FjsSO0TrkaoZawnZiVV+DC7R7jz2AdR7phhhwhw7suyp5c5CckQ37Di0nMWQlyKBYs
TKXI8f4nqOwOCdEwhOBhNn7JbkWrCduHCgIV0iv35Jd0jFVPUmhcCbJKhpXtMagWykp4QPQl/+yA
fZTxd6H7LiCIitv8qWzpcN7I3EWfVEmEKBMu/XFUrfUX24RZAX1S3UAqqD2kjycxmC/ip5j8hP0G
TPKHv1S4/HCAqF37PmY5UYg2Liop/sv41OmaE1BBAqnK1+VFBAG07iEdERuxEi60fr14qVrT92Rf
tNenFOkuwKG0yun5Sl+VVFSvtJq60fWVPRTuiPYkpU+v58roIkoBwclPXckCzGEwq9XvWqRoJ6Je
PZEhEpgrdyY+zU6hTuUvNaavvd5Aw/Mmv0z8zN6bcuRDLStc6UZIFLKOvW8Cwc5Gd8/fgGvXqRcR
/UOVbMFDBq3Hz/QJztn4Q+UV7+SNpx/q3yozD47xARe7uq1araKz/tUBmAzhrqgVNBkOeXbxfkUG
mU0zAPG5vG+O9efZc2fbqQVKQZfh5g+UL9sVydOnN2ppXj5ZbeJzU561MEot/+ePQ7D5Dqwp7Myv
VUxBj++MJrLh+FWzaNEE29pjm73eJQiijixowe+51vXCJEaJLGReXdfV93tgr02Vv4FAGen+uG/i
mivJoZAPQE4Y4DQ3SZm5w1slY7zHuTuPdE9gTuj9D4cVM4BRGKFlwAu76Ic8RbZEQ81o2S9/bG2A
KLGY4QpBUUomBmpfEpKC2SAIan/rjFL28G7B2Sn037OJ6hzVcdOhBYYTmGBBbOROL8/PZRo6f5/m
hLcXaOuYiCxdsnydLRPJooPZA8DD2fe61ofeQU9KgfFOYGH9N9KaMXad5Tvo1fJIMHtTQRNV6hNt
W3BPNTyr1jLIE4yW/PSobixIblgLyE8lguwImGIgJD6TNGMDDLCjRVDkchNuZYl5m6cTiBlaqvcE
wMGXwjk/XmPsWFJYGVvFahXLyNr8GeIzPnCr9v5B6N4iBNB0/sNNvPWtcgfwCHDrgHfSrBJYIuzh
G1Jdr44ii73O6jgnkKPRR+4h+aqAsUpldP9W3uG8biLMXLEUAc8kmV6htPX/Kaj1c64Ny42cLlPj
QqVI1nvhcls/H7V5fAP4I2yVbclKf1g0jJ2yUmN/wEysUyxOExX9IrSZXvq6wI+fsCgMyQtXfwk5
78AnNfFZTr+na8KpX+OgsvOIuktBaFo3i6QFBMLJuN23ght3Rp12UIUT7K6Hie4ejFDvd5C5JCx/
g8Diks88CcCXDi4qfHARuDxiiToRB8CFbMnSAMx5pZQd3erEalYtbWd41j6Ka5krtAFKkx228Zdw
DGe++crQ2/q00AzVltYz7EttC6RUqjRx5rNsRTk0LYYOKYe8vnlebs1nPGjE5lGrDDqjTkdx0lII
NoPtG13pbSi7UsCbWigrEsRwsyrmS7xeslJBp2n1r8dpifeFz7pc8D61CA3ocNNsuC3Ct9B8hEb9
SSHi6EQgAe/07ZGjrepONSsnIaZOt+CayxEx79nTQnN62oQxLCbPofK5sIMtPscHdWGmZsT/AIZa
R5IVdsSL+zzwgq6bR6NLzzfAnVR2G9ziXUyxnsowYDMyzdqQvGxu/bgblPdoOyEalDGsAqlvEVyV
CMxdpenVROwuOK6rB54pjvPxwxTsfpCVqcnt9p9zwiKXucnHXLfl70QPunIKVQBzyTVDVxb5Qrci
CocqyceTRc5ji4MAFsx6mOL0qgrNgT6CXaDZJUH5/z9oLYdWyQa6+ZmGMuwKrWqZkrvRKGYkly12
v3JHZPJiKgTfZ9CqTA66BgUY2DRRUZXhS+oZCtB+z209HjGMjYy3fsGwk7ovcuav/mBu3G342xps
UNzEVuQPYDs8LPV/5LZklIU2Cv9f0o28Qjqp9KZd3btDkXMYa+pJU+ShUk9EQf7s8m5ChEFxgZ6+
EaauEymKsnT+ARJOVkEBnZlhUb3ZW3hjHL3v0ENXqr857sz7QspZIJ22bhwZ5689BBneTURDRvIL
0AU7W/KZNsWQWeRBUAn+PWXDVexb1Hpc6kxAsH4oPJjzR9mR7riYTjJQwlBS3S3Ki1G7tz56T+O7
FjFUcWgJbtXPmyajUbAV1u+Dt0YlezPVHG2COG1Ksc1dsjwO2kBSvA+x+PC//6ORsbQiCz/Y/wv+
04cG4zDMuE1zJ/lP7cahWcl+DuZ9kGOBscT8l9EvYazZmD6G43qPibFwJr/hEgFwubVgbikvkZ4P
Mt/ENcIqpnzp+guj4USYEsFNYrk3PY1joEDrJJhIrRz64h+fnyEb4uFGyDtJJNfZKHlYza4QEEOf
y8qeRP+quIsqgjtcLxUtvIFcjXcs9NrxxVgPG7/V2TYpRDkbgF0fMD3LWzMw2vZ8M0MvbB3DdpSH
du8UuuJNnOe8Q7KVVckMyLtq28MakrIEPNl4MYhXadJ+BYmX1Plyng/j7EalOUTrAQ6WObqykpTu
/AxdoNK5tjrhzZXgCJwO32NsWh8cvxCOyB+KqrklWiGOO5k5OCpv427vbJvf8C5iTjmTanSA2ziA
1UD0ZKqt0x2kvgxzLa4riUTtb2r4hJf36CONALHrkihhJD8UkEZiu9TORHKpo278ymm+RakxXg6Y
vLFJGbkXHrJovc2zMSCTRvL8Bv4M5bfBUuOGkJ3WRSFtgDhhO7LOrzgx+pKMbBhUqBSFQLsKEtYj
a5WRGREMpXhj6tFPW2npOutxhfF/i9zHTLuD2/mnYpXXPSRUOEki8H1uXLbQZGaqIsV1S917N9x8
zdswfTTgiU1moPo+9UM5e8Qtrg0VPyTfimg+q2/tIOGO972GzSps8avZG93pSq4FOTfd0B+PEdHM
Lg025aPyMBkH09Q3gcg1ZvudngXssRw78FohF4sQVgZXT9rGf6szJWoFic2DRdpZTu8FOvkmTUva
o5j2eyvkG+D9LpIpA5TZCbQtjkValWMFRTmvcOZfYgf/zaf/ohafS5SlfkVmAqyzpjCSEinvq1A2
yHg5BrN+J+OEtCLi98+lEnLagNmta8vQbqIR4wOT50PrXJIpHOTw4WOScqXSF84K2BPYO2JASIr/
D8HyH7pQDVn4rQsYQAs2/9tUvHVetKNq5/RS7W/Y8iONFGzRmFSXAtVhgT2kv0QpRzeLGvi8oCTX
rppUInX9bL5dlvsaYWIAkcR63FcjUVdcJBPvr3WuBwZyY005D48Vzd/oJdd0CrEgujUB71Ocg195
2cQ0XQvTjnmVUf2Z6GR3z4N0L5+0molsVuQfaUvTDNBV+kqZ8Xktv1QNFfQO+l4TjlqN+rrVrRvS
s9o+wt2M4h7y3dLuIhhCYskAq5EP7ovLXq9E2PVpPB8PDQmWNFSmd/ukOcAX45aOnp74+38w81r/
O2U9CGUX8/B85aQA+T997Csb/HM6+QLRcnr8fnHn5zZcWeDwr7NrrleYY9c6Lu78mHXhY4dm4rtF
tHfZYIJdqehAJ7vub9MFwjeb33Und39bqFEpkYk8Hw0+vg2HX2YMxz01GiWQivfrv4OMPIq1w1Fs
49S5L0ck1uUex8XiH/lxOLelCxPA/ww5Mj2YuvoKqHF/CCtQx+cYvJ+lT72brjUQIzpoUzFLFW+c
3MqjXP5dWiZQEDulLnzCIn9Sd+69n0EMUFcCc+N/Tc5wIwBjPIC55VFmGTDeOfPwo+vUrR67h2z4
rItpmPAOtXeMwf/Kfntl1ZWn3ee7BdM+GLxmwPQAtyk2Otl+uQuYcK2hPoc/teco7CL5IJsvV1FS
g0XjGUZIt2051cdXNBEpOUlv6N2YWIEp62xvyR6Zqc/4mG6wFtv6CquWnPZW01hf36TtR/RzbWNG
9j7Urt2uIgjhjr5XYxQp5gBg5XKLlU3uLFaV8lMQ2EKuf2solc8kCVU+odGff09S1CbkVGWpg9GZ
ANGMz+yLk4mLW6eQbJ5OhZKDvfypPjAdrR6d8iNMgj+DIIxPJTBmnMnPWvYKELwWZOlmg8i8NShG
tmIwNH9BJiyVNnrX64+SylJvv9lVHWtQgAQL+ekw3cShf3cvZlLae3mVuxO95qoZAbakS/zwcON0
2kvUdnNkUnBshTG4NtSQdQLjekOXcdyrfhdBiKN4yhF4knM9mKSc6CL8HNChJXc6Jsls7DSLbbL7
PXjz9ajP4Ja7oWm8GFuu+LBYX0LcBXWwjEhSN+VoVGvHHbNiptcyP2dZ16gV1zIBd3nZnCKcCYBM
PyVEXA78tbs/1StQ2gk2ncMCrX+OGTZjvlpkzF32aB48QrvnsKV6asYV7qb2FlUt5Cu/nlEuI6Sl
fYF8+d81ZI3gb2ZEnGd5jwI7964m3zcVwxhfVA8Cpels9SNlIUKglCA+E4622pM9bWbCDbA030nB
01gLJZIUDQ2/6celqWh6MHl4Wq1d4QjCIic8EwnqoutQKfJQr4c6HyJqb19UhbNVSyq7okDOq19P
Su5W+BJNtWrYrQr317vVWlvZEy2fI/MMlYvKmy6Sp+DQ4MVPObbKnt0H2cgcUDOqwFoP6xDI2zuy
Rj2wf2UcOmdRamwUhF5rwVFIoBuiJzL+PkozAguDAH7MqHqn9YLAf8u+lp2ccRxjOTZgtzhM4dml
c9D8aDSYpFep85fPp6jRKryby2ShM1bhQhEU8P7n3svOF9FKXYfMTQM3NDcw0HZqdZMWplcLcL3V
jxVDCqMi6o5hUcbOK6zR+sXqoU9F+sCMEnCkL+68NzzYDgMXJLiQpgRWgg10cvYoY56b0fpdpIEg
IV4W/Qnoqa5bRBuZhdtO3B7lVh/5zWRd6SE9jYWq+79ydSsZObfs0osUXPFFDxHW0LA1o3KWHuLZ
HWmpOrqhyVsIEVuQ8TRZ1mxQ8FVx1Czj0RN6/iDMXkJESqhcWQSwApzIS7gEjbNnZOW1fN4sdtBU
lqhmP6NKwNXZldOyUzyecRAjz/TEO8yl+JDAGIJVvYKepFOUXNJlC1XGbE6Zqmwfik1NiOSzJ2jz
37/Ui4aw2h36hwNPUamC/csAN+K5zb6aifcg+ZbQIklpBCWdOlXbGcBNw8tdxqWhoep56sZBFLzL
fy7fW30mbtIyod/uIMDrNN2oAV/vkX0WXNd5MGtCbwsWXaJbxcO/NV7RbEr0doiS8FQw+Y1WfiaQ
E20IkIlOZSnFrV8luAOavT7zlrHvDjz2Coq8NWgo502zQ19XfyQXnbCX24SToGpbSK6xy2HeyfQk
zD8kAHlGyyWt5Ocp/HStMJjIG3f7b9PlfnY4PLa2YYjzeJU8YnXpKV5L6xbwck+Sm31kIB4IvE6H
cjxmbAc3YEbhe6yEurfAA9mZiTpqXipR1VwYlGj7e/ru/TLlU6vRD+QEyDYTF71femuPznN14MrY
5WillU0F9Dh5J0vH9jJpgFGMP6ZgxWQxV9hWlUeD2ETUnv6SkqjsaTr7w/sQBtXzFq3Ari02BFX3
LAPWCU102TGhtvXo6hWpZwvcGY5st+Rh+JcgYImzQ6OKQEURP5VM5n9WBSZkixjLuZsqK4YinWfB
Z9bXeg24JzYYBz9leLEkMl6C0oZbhfWvt+qAstEBKZV3xASLpBRna927LYdWPPE6sP5XY45psvUh
mUBYkmpHGjdpfPkP1PXaWhUzBVeVdHwm0C+fSe5FKa2+gf4oECPO/gwW3dYE0o84GKIBuNGXYXQw
gxt7sew18M01c1Op2FCJXjEZH3XAS8pwrrZskppZhk442GNNzPGWTjfMgifs4krUrCY73K5HhQLm
cI6Y9vExRQncz5GeO3+0bKufiRQzG8yUxlCZWMYZmg8xJCtykxhHKChaRP4NFE4FRJOG00X34f/b
a4MeqysvuY0tbCsn4zVkfN44uF++Kzn7yOdAoRRBt0rrsWfiIgNRec7zu9XLd/fnOAyI83ZOyYlg
YamYbpjoXcLOUb89ur2DklTDgJiDovp7hay1qYwoBKTyqgk6NJOI2L5o4DP1y0H2Ex5AWxEMj0dS
6zczL9al4ZcgkJVnQ1X8wxEe8utI4PTIfj8UyJVto6EQea7O9953XhDw7ed9S1GTXRTPcY+ZtxQ4
1we4v8ZcqDbeSDFHqtC79miuSS5DsZ+qrhyj4Do6t1pluKfXIfs0PYnobFsR8gG7mJjipyvwv0LG
pxb2hHhdKFjNNtTI8d1OpSkNE3UBQWKmp+0JD/UpdCBEH4RrTHLkZhStY39RsiMFhiIViHL6U1P4
mu8tC4v/qx4XlvcClV+x3jv7ykp1EG0Ty1Q5HKGPao+wd78seCKCpiWPw3CLUWa/NN0HHREJiQEz
XT+xQdn6RtKf3+y/qYyTIellIkdIGJVo6eCqbRJASw9bnfOsI6E2i4EvDFRHNx3ltw25/QGgupyr
eWX7b41VoEKcNI8VaeulIwZJlIoL/b+4WvmBevRfnGbVEStc74mVOaui35ZkZqykEhr0GHCSJU7O
w50V6HpL9t11FkyNzOCD21XzvUVRPaEERZ/0EE0oCSx7XYJZ5E1t8B+EjbRIZ9sHP6ds8rhH/hlk
mkiDzvwIW/UysVi3LPEypGGCX+yypb7WLoZcURNMAbEqZ6DFPIp9Ypqs7OmEiwjf/PtieFSMMTVq
Q5hoDukEWxDDGQ1qD+5fP/HvyJCFhWDcet1N0j3KBjIpOXaS4Ql8G+6DVTiRaHu6ct3KEJ/LK6Me
8dlFwsl3ySd+wryqIL9W7Rd3vRKwYcjGk/+NuJ2L/wSg4cdAFQCCkAMsQxGotN74cH+jR6PqzwgQ
1AVL2eHLXcitoPVhZ01MY2kqGOqJ0b1aPZj7TkxCyHkaoIcuklkeas0WKrLFc9X+N5r0C7IjICgJ
eSSfQlrcWefWr/fyzXD0KaKFQr0ZftHEnOovaXhwd7RH35fwJjLAGMaRdtQB68D9L5/cNPJNYHIe
7BWNLB23f1U7FxP9MIRgMlm2KEA8bMR5YuIuVLoKMssBeljsPlZj3CjG66u8cpFhNrJagRKNWHsx
e6qN3DoHaydG19ISykfE5ktrfqZ5tIO5l2X7jkrdYWCReMIz2qeHbC0Z1u9TPO6d/+uD0g7V431O
xGis6pL46j8dIM8V7ioH3jBOXyGTrWzDbv2ccFLT35eynqcGYv94sqkOHB5mU3rFyda43bnj4ZX/
dbRDm8Dl6WQXiq9BPhKL087lhoc96L8YUn/Q9dgPDC3blRwUQ5KCTfkmwaetHfTIlVoEA7S91GJg
gtvD9uMBVaQCq9J+lu56tddfVnR5XXwlnr/YQw+vf0PVLLthEk28/vevFGTHbRVDTbefBtv7GTsf
mkP8Ty3JR+FshNcQpB5r0pvnt3alxT2k/oRO1k3B0cdZzxkCaEGufa1FB3sufXbW2AuvwQ64GdjQ
lIa6cxv/2rWGMEcyW50bgYB/fZvzGAmULazPB/UBgjjDnWgOcfQqWllhNjFCxRmiq9B4tM8ejZnP
5r8BvKzZEBpsCFFjWT+hpWhJvGN3Qtc//F/XzKBZvuUMA9e7S2P8zkeBKdsW05BEWkir/wsqNeYd
92Mh8j2/DAWNm0gFa87rg9CUpJLbvCMusgGynDr9JG8ym3TGKITCCgJ3vC2I2cRTLs67GT6+vM/E
GWV8J/l1s/qWfYRbaThwfg9Nxjm1IXS6uh60Sw8qGhfKB1RnHrjQIGqP00d2g9/AxPkhfO94gumE
II8T4vNrrrgVJjtVvQbvZgZvGiHjANlix2i8H6C3Zj7RpF2NtiPPAetTMyt22fkeW14KVAdNmecs
7ErLkaZAG5Uu1N2TxkpT2JisyQDIAJFUknx8NyX/wbemJjWlo9XC+iIKCs8kWQ+EIs98V9tCgMBh
lmLBXmEcmeTBrN2T1e1ZO7LGZewifp5y17PAGKJsyv9LvNjjcpvTExVVoFAM9BXf9ZP23FLHW2CB
qup3/c6wBbF0NGfgaijpW6pvtlncs89UUgAG4PONVW8E2+tzK0ZBDQpQ4/a7EPXPG5kPSOUYEI1m
DueRkzf2F+P3tdz19DcB6IsIm2ekvKp13kOE9dLEleBB2DSyrPsMA920k6R6kPvl30gmYu/3KAxR
HBfRmWBUCk6XVNjdxLzWsdp5SozYkrH6LxAHvVH1QKgo7E5b2eRLM5wh/RzxTOo/ftTg52I5m2Vk
l08IGnvu1eXJXqwC7yGuoL6drqmSZOi18HU+rkzpuvVdSa3mM4KMGIG9xhBUbi0DCUftVC+ImiZI
tosJGpTshQpGb8RkN04pRhI+b96Bq78MDZvzI+Q7P4uJ3ujXyOb2tSz2NKmIHugF+n0nb7HDO13d
TC7n0CKVlbBofKelVvsILFr4ikUgWu1CZwT2vBUfiskzuVB3Nc3RxFWkKsUllZgKlvOn4Ztr87K/
CLnAYn9y+ntpNUBtIW5ZV3OAZx+madV650FvU8hb3dDsMPV+1QRRPB2o5gwMbmCShPnyc+X/TWzl
PWxm7xL1qWdFPBfck7TlSdsQrXxgZ2V5taZ7YQzviEoMws+lfBTr5sTmfFzw0dsQyVqKVRjPKFE6
Ffpe3pLlJ1eKYpDS6SCsCC8iA8vMtYJ2cyV6H29F4bQYXEjDROJ7cxAwU7ar3FYhqJ5Z3Aec8+/c
fTn/LfuCyD7JO7ccsdNf+Or1BrgMZuKCxdiRMUmyU7wXq4i7rxMuQwlLb4tD9mynvTjXbAnMYV6P
o0fZpt8qe3l/lyBj6wWyCIg0yrE9F5ydd8gJTnu2OouBsukcfNtZon6I/5xr52NHQ7iS7/wXKcr0
y6SvhZZH3kdK+PozWYFmkfhdSpW3e0TPzdYZHTm3LZOUGwYXD2Z7Ep+LmFt4u6YQ/07ZqF9kh3qn
H9WF4jrmJVit5h61IXFusliOramBQkRDL80QCwDwvKPQr92brhjpfVHmNl+XTbKicPW4YqDmQZwx
dzGv17P+JbBro9MCOyD5P5ZXqZ4+0kdshOFKcw4yONYv/M/DAcBw8+kS3WDFAdszPgUExI6gMCwT
6zMPMaKkl4Pa8Two6X5gy3AK2iyAQCIEzXzLVW+kYl7vAU3rLC8Ip8keiVpbu2OWPmB7dOT3BAp3
WQgR5puuin9w3PL/7eSwSj2LJqorROqdywwmWIY/tIklG5n2w6dER/S0fm9f4144HvJq3sEUgmXj
Yc9T4v0/G79TxXB7wUNrxN+pEsEbmFrGYdxywK7gjUrZfuhyPtb/A1qb1XvjtvPQKi+IcFbCBJ7o
C16sTZjq7ijP9ODFXBfOpQXq6sfJc+eD18KqdtvUbL+l4YeX7QKH1U6UlsMQj3lV2DzzoCGI9kvb
fVAuJCoDerafyJYold/ayUbT2m7XgkwpaWvoeYR9OzP4m3C12UVRU+3xLV1nghUuC4c/VVWNmy38
pQzaMhgrvlub7ZSTyUl9RrQovBETdXmU+h6Nz/Q776queadevMXF5RNVF+4szJ2aM1VmNIKzLcyF
LOq9bkx8UuUsrnRO5ICE+I2eTfoekAoLRHTHMTGbYXNB9XuOKebvgMOM4Vb4yrBWedjZZG0Khk4q
EDfzX4JxTn3AeJusyFUsTn6XRWDTHj5otK/CyRB4aex1Mb68OLsr8viIYbkpHsLok9bcSZmXwt8p
WdKyfrMeC8xduOdWaLf/B0YuotSbBC6iMWcO6ju1Rxm2PdWTSBGpHZYqYoUbiAGUZNJoH4C9FtkZ
c+FsF4EwKXdImXHu691lntTxRXYjJ2Hn5iD44dH1HC/xJqAEsC0T8SOJdpBLTnXaXXqL0yp5KZmm
wUJlJsm3DM7O6/H5EiVKAQx0FviUGkIFULxZhh4eJQDoH/4eb4r3Y3RJn13SDTm2yIgZfMiWKo2i
+KbbJ+/HB+f4fuvyxsdwX0XoGTdzjDZ68ywGjeXPAOc0+tuuJnpW/GrczxvW/Vmc0Kydn1+JaNhu
Sa1hx5b+CXCVUJFj5WMpaEkn21crAPU7nvHE3trjERHza8d4hRpVeppPxq4/RA+iJCl9wr7k/SZE
SxUhqS8I/96DHPMoMjVPaqD1wPwBzG5mMg1Dhqpgj1v9Qjjv5r4ig/W1NYmiOzHy0CqVzdiq/wU0
n/KGhvg+zYTeLzY7lTt11qhInx5Hg0eEua8S7O/ixNXGtKHpKug5HQpAird79LjprHvC1Sxkia1K
Qm9T8lbjhfOuaMTkzXx7vrZxixyeF/c=
`protect end_protected
