// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
lUuYxnQsjbb5wKQ2Qn3qRnYDCv4wLVbpU1i2y+y9b6jA8tWje0OUfVNqpMdEgelwh86UQHehKMh9
lsfAIzCdqzfoQvOu9CWn6/QPtfi3Frl5R28TTPZsdbVKxd3oyyFnE5+GMDC8316UJvMBystJHg8L
kBVIeSXt25AwLoMVVtxMXqdBpHvgOtJSbBLqAdg6WGwClA6dTmC0eIplmHF6aDoaWhOJJUkWdGpL
vDopsmqNdOPYDPeqDLhJNww854da+ndft4V/wKcxTusk/KtGRExbdjGmv1fp3eGdHvqnqGL6oMXM
dlT5NrfkvKGGkqn9wfDDff98Uytn6PzA1tsgUA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11120)
LEqEYyGi4H3dw3xTFyANdz1Tw+EN0p9ZS+Jrd0+r3nXHxn0FIjIhifh2SBPhQ2nFXzQMFAPwgTGg
ZHhtVEDe9Vhwewp/W+AGT7ZAmnVI2DKQdT1okNB9lB8Wvcv3n0m9SSKx9qns2RinTmJnj9f51LoA
WjLNPXojM5RWYLEf+eG/E5NscDeIx3iuo7Gam8SLk9opK06xfCmFh2tWY8VRAbKu9MnH2NcwVh/b
03MajxhB7K+ur/xU6IdmiaEcw7WUYMc/3sUv462NpLny9bUbL6beuNeMMrUvMOI8g2lxf5YuV2k1
3kV6zTTD51XWilHg9Vn7tu1Rvxd1QCUw6BGANuutrpQ2+u08dIJzzbhlA9lHWjwS/i5/7TYCZrk6
JCt13XZhiuKnGV/EfMeOB62tQMwCt5mAaGETGDgsseEhn4G3aycvvBN4duVkxQCnBtoOVjWkAPbg
pETQT4tLpl4mdkYwYwlTA9q/5SXNVi/zMwmm/fpJOeO1neZ8s08GlinNYD/tAEqI7cF+YNlEVr4a
j+c7h4pcpvobyrlgHxfObq40f+rclgamAENSsPyDp28keJQsuVOmurnzDTSY2uZeemcv7K0gqpIH
QMcN76r5i5k1GHxGVAiufnnhNKFGnlNT4SAGtMZxx3bso2e0+ZexZpOy32S/41BVYZnTnLl6UTYn
C7fzPxlYE+mLj2EbbHQuwbTLNqUeb09OQb+8u9qlvF7BN+E6EZkBwHf8GbKZ4/2XxfurIvZZcwxs
rfD6iQYsf4tCsdYWnWnfrhtRSYWojMIHjkjnL3pc7/HGF2VaFOQtMzWZTFmfN+m+a7P8exwRF3q4
kLJgjf1tvVJGfhxIueVpFeXMvDOmJm98o8z1BhrA//+JfceQRsnbcdJMy1iACg8bTrqT/3r+LOtR
Cc1V2rrkQcZhDx7pSvtrWuRwqZrlp9hN6e+cANJPmYBR0UEe4NYQ1326Abao4epxVeBMllKq3kgc
JGOba0GrgMWqp6yAL1GqDPwDaN6LwUbqo3cZfxHS4QjKFZNR7tPtPkZn6ylpqS2qZAMopx9hl/hY
wLIB83dIjt9ieXRBNNosvPr4sD+KEKulzmM1jdf/jZcitYHW39DKSeWi7I9yZVgREFgUZB6T7iRx
uYHjWFf28RVkAkbTKGeQA+o4Y3vLL8NS+zpOwofdMdqRJWMdvJGrGzBbM6k2Kooe4dlVkmmXG9MF
LLC6a/J5ssK2sMxd21ngyfFgxKUQXHTTuXEDsW3O+gMRhlxTv97X5SkPngvN+l/jG3MMwX5SB0RT
9tBsATstW+si+5mG0PXg5CEj8MV0pf5IzeQe8p3Y2MEkciW6FI/2VbKuyuOaSIzfZiGuIZx9IyAw
7I1qMEp2YM81Av1TAZBoY1LUm8iejqAy/W4kLOCbFO9ceiNKwl5XGLRNvBZXYDu0uNMX3E2nsAwu
0LnGPw13VGSEpRFJTrTbhY4WRuc5xwo19Fv0TxXpWlUIe0OrQ+4YWGaN6vDV5pVIAOxttACKwV6F
YleJ17noprkZlD3haTi7h135SHs/6mMAGtZyjo1MBYAZtI1IVEZjSKFMVudulb80B/VfLJasfy8F
zUwnXooAQnm3tO8jgpuBYECMrMKjIC7y1PKPia3tovkLRvc9pUz0FMiv0G7OxH8hkOSNjPokvJtx
DEcKkvXczilbjznTScuxcSKBaK40ldOrByZ81UEW9coaGcZQRWMMNSqB7l9CTKSqI+cVUAdj5i2c
y3kB7U5VA25oGGM4+FMOz1xx0narxB5BErGAqNroGVAwFvZW5O5Z+qC0Yf+WYYkFezdG/VAF2B0P
TCIT78b+0wsWoVQMjxF8KE8WsVZplOpL0xJAdURZE/wYGaIynFmICld9wDLUl/9gowciqkmIIGnS
el4feTEDHFdI+A9hSbAyzU5kvZZLOj7akxB7+yl3g5uxm/swM4djDykUJQfS09wZLSBsAtc+fODr
x5F9e8PycFigO3TW24J7Ry3NyGswn/XnJA9qidOGEn9CRXjj1DEXG2FZOUt0lPhS7UaltXZuSU/k
pbqkacxh2zjYBxX2uzOkaH6FF6k02s5QSsQ3n8MLpoE+eNVvcNJ9gYxZDVSbebOucY1XBn7/CP5g
IH1kHIQRyV9pdpgUlWy7TneoBvypppr9WrYZm9u6wLczDOLwxRgQz6oSUMrggKWgB5P0rSB5j0Wy
I9iXK/s/yCMlnxxbj/vSqRkprr+UOnIelArw9g3UcRdWttLh+N1phixltEmvSFRj0fXK+HMu+6gB
559OG5ICXxQ2cvQBUcLEAaWLj7ulKP7y/sGc5QqRF7tPuZFtZxaoZA/PwVsjFzgxfRr/9bigBYKn
N/aRaKui1P1uKcljxj2j0FEmn1HnBtYNjkSsieh0o2SEFnpjqcLz9XJLYYfol3VQQbIykYkxp25X
9aNBamxDVkGBtwHw2p8U+vCyC4cdUSDIcsdbXCyYloCnHN/x4YZZKc1y32COadXFDsH4pIwNt/y+
M1D6q8e3M06AvEW89FjM6l/EkoXFe3FiDhCxwbmIaTP9fS6yJOpTZ/3Uh1NYrTvy0WK5kVKzYGuV
PC4R5Q5SogyO6dcZh/Dhf2J3d+nMwUi9HNOi7ug9cYT7NKXImBMMR8pdkUUJvX6CLL73ZwsLgV8E
fH3OBhslQ/GD9fyzOEgYRWDGtsX/k4llWCNkdw11uzD4K4d/WBLMiMOkRDYfPP89PsQtOKBoyqbb
ddA/XiQJOW2NZ7f99oF8+3SgEjd6E3Q8PMRULTVluLEw15XqAih/3N0MgIPov8JQ7KrNS35cVzMy
G3xqeV0WDUoh/a+S+8s3y7RWdtPtTvElz/wA+LDffEM8EM5WPbfmhDS7oq7NVo+R6IXczsG3OYsn
g3j06DPeyxmczd7vWhDKsdhsa1yx+Rf8xBxwU/9M4Pw070y3FYwlDPadDPqkZ3iaCobR6rnpjsj3
Yc2Sx+pkqG0YsrKAIKTjwfpwTXflFPK/BlEnlbOcm6/wIaAYolSkKfa/OBcswLCaXue4gihfy8A1
qlYwQTxkSW8/LdrupEcL7+dbb3QHuKHml5bMQ5g/wmUY66f94vd3efj1gWyUqye+kL1BLuKfFRTt
mCiZ2U8rjrxUfSUGnKa4d6VCse9k8pQLoAaEbgm+5c6ognw+Q7xUowQn+5IMvpA/TuTd9shyR+7A
rNPzdFGXThODaPqYSaxBBpJFjEjYvJQ7cKUpN5o5p5w4MDJj8dGzAKEp99VZRzjg//y6Ziy0L8vv
DBiF7e+qMcoKkUWbt60wEoAn7H+h46i1+GbC0B3PAloYrweDzCieskQtOnBJHHZZRJsSsYDQBdfR
pfmzPFudlWjDCpkbNASNa/1/0eehwoGlXCOTaYiMtNoJ9e/Blhn+PkfFTJfc03s36AjIQSWl9TbC
+5grONyjaPb3EMCOLLnJV2Z3fseJ5NvsOHjCCoH6wCRjr9KAus1Ai263dn/3Cc+7Ui27ThmKkN+G
PDr4fSaPRuknfpFrNw9NeGsniUzf+3QuDSLHwjirEQ/NcRIMouIL9ePwyZU5LbaE2pkffLglSVpJ
K5wOvLGkCS/p8796K3J0H/szZoik3o7ZVCvboml2OZGoO7ObZpvtADgOQ/OV/HGLUdQ4fATCSrSf
1vBMyPLmg7wod+yoFfDdPfP+EwqTCu7I81YProd2XwCuuaguD2FsUwxobE5BPQ7/fl8VfZ0gxno2
5R4/tVg+9OuzRXLgL5qTI964RsmyM992jL/bn7pFglzw0m9T5W3cQLjxgIITWdLZ8pUVrao1+qN8
R705rxxqawpPgo3Q/YQsha3zbME3zx92bdSc+TsZ6UeoDMTEBcWuZKwMG+qtF+4r5CpbpJkBgUeL
oBcdc5QZN6d+VMPoDbNTO5zeydXSPwAMl6QVBrnWmzSaKUJ+NXAxjw+vbjJ45JYenRAAlvq5BPV0
7NVam8R8JHQDl0VUXrYeq6G1Eu4x11bU05XhxZ2FuriYLQ/1ltAsJ7RUKCKexvCiVTGsHkaIKs+z
jOsRTl4riOJ4RnOHrN4uC9I+B8xKhU4ULnAHiwrqgW+i4UlcL7wgIaRGLBH0STnM3jzQabxzF72m
zXDjhZXtvhzpQzV0U7QSM0qQq6ZeeDiXxkLGVDn29xpFWwHccxyeSE29JmD5h1GUOfj0EN8NLlBM
9EBEfXAqfDK5wcSRfD1NTpdfEy3vpCZ9bve5CM0ooJB1XYHIVH4t/9qTFqxszn18qo+Bq9xVke5l
awIiYRHxZHPg8rpVHvZvcF2f4V3O8Di+JKhwfNE9TU5/b7ICC/WDK4quDtagWF3/ANx2Axvu6ptk
xMKYG9FGZ+g5zzVDLe8+aGBDnc1BL9HXJ121HUftoVll0qVdG/mpg/xrkK1DAiKjfnVf1qmFdvsZ
ICBfudPyTNgwapijsEs9D10N+jvqIWC/HyUxS/LSvqBRzQIt1son/BNtuvBjuCzBYZaA0lmbqtAG
EVIvQ8SrAuYgxD/k1zP+egK1X+wvXkWJqr3ZgVjM2twbsniIM4T+rcSSiS/aHGb1pe+G/iAeV44k
7KMDaMdjGyr/rHe+C0HIAoehR8/VrEft5opPsGseWiS/Yy241OQH46hHnXceSq7lK0q01oOQjN8k
kKGFFVp1q7c33BN39zoHrpMFYFx0x2xrzxkxDQjeIDAlzAyv+Cq3YOEhyEr9Nik7stOBfhIX2Rvj
i3DmYKHr0MRDR+ZmIFrzZQQHrIP6Po/Dtgw5Hd/pQG2g/HMll5bR09yHnYTPOZoz2Zk2STHbqZIA
Uf0nb2VmFt5M0GBOKLDPQFQQBCQ8YxqCuapgwQ5fGq98jtATQpieB3spOp9tdLqlbKOZLQCA8JrR
sswhZ7nYRa49CVcoJqFCvgPNz1nURq+ZCoAWVHMtfiq5DZU54SbuJUK2frAPt6sWhJKnkvVqQyFz
mLN1UOQ/r7sh/oe++s2svk071ALi87B1NKVO93PPsY8qc46BMkPg333kg/CgpXrAshAQc9u/pMav
+S5hSnyjk278lcFrCU0GzdGaghIOJREzVQhuooJ4REhPU7mEhz1mtXVuACiSfbcVx0dFnsapWpmS
i4kdQcnvbP06tK+1jtiRAXGrsMIgmmCOQG2ZLOEH3eSAUhB/PZ+8AwoyXlmIdIxjOf82gU4UrwuD
ghgIgZamBJEcXnPz0nhxJw4Gzq8LIBPatnT15dxuVjhnAbi6BJrZuvT8yR/IE1g2aXOkjleTt4dZ
tozjJiBdSgurlPwv9AAnlCTSNcZ21Kgs91bEWgvTcYgdMcms07kjB64ObtEZDJ6/elhGQbr8qQ1s
psplbKdl7cih1eeHnTmVRpl0isnW5J03pmdkhZ4Or93RnXHabPspgmCmKgegqXoKN2oa8JFEnuiu
apRgr/9jaSoSKcqDU6qNhEvXvc2syrC651NM6QAXNQVRzsStt8bJ9oYF+yFnzeCiosL1kP8t+xNu
2X7ki+cFWQMdmcZ/sGs8MoPMlO/ruwET1EeBvsQ405h0B+CXUhAEICMbllIFhUi0gMCKvBY1pyVj
NZKotjt8d7NnRhpzt78OJyxDOIMATekzTMYqFAULAww77IO/wC+HYaO8liOf7nREckJC2AF6NCzn
XML/Sc3AYyIUCPkA0lGVA/qZO3PkMYWX93a8cXtgbxS1EAupKHuQamwFVyzt/GGOsc9rSip/CqmZ
UEzp2/DXMMYthYmVPkiY3oKWxYGsjaP85f/5tDOjesov7QaO3TQDwuu8+4icXj61tgXdf8aTY86H
5+cqIqBu28SmbHm+aftoNNLppkLJK9j2tJG+dWhC5A5JU2KiVPqo+YWstPHhNI31w1nHt8JFxZyD
7E57q7G2+5kNWr3YQT0t6qg8Aqs2uhCH1GdwfLaIwpJPo5YKA7xq5GjFvMarcUOzRemuo9bMX0Zk
1k9iwkD1Vlk9rO6Au42NurUTyTT4dkDmt22Op0GRoVus5IM/7nAvhHXEJ2Y/rBl+IK+ihQZqL7Vc
gF+1ZzkalqNI0BKuMfXy4p4nWpuPWwvAzAAju73Y4iidaaqFm9hG2/oZfiqUa1/Sir5SNVufkfcS
5vtS7UjWxH7kXLOzbXMK69/NmD2hUnCekeKb/buNxq7JKnRsAR9U+Ap8j0/nPHs3OkvsdX9UB6aI
xZplpk4oPZy/RIospYBBpcZhGWE22XUsU1EI14dyED7+iKKWj4MU4KLMqJSQBBYltn1MrmhaWgBB
1Oxg2S+USu+uhrDsq2SvvnOLKEtdUx8GRBVcHBIP9OKvdheXzF43etCtsQ4PoSIprdAlbOM0DkWl
xU1RiI2RhDsY1aQFJ/iIjXZ9hmwutmEzYW+ExqSxm0LmhbHjBtpiKGinABEsEuZ1+DZlGHX0fL7i
piSGeUpjET5DuAhF2RA/Xz47W3yrCQAtQIzGJMgwXTGHiXtO4pAMGeu54ZFASa6XoBu1hDn/gs18
UAq5x7pJUkf8jJa0TAt1okwvcaWcQs6mO2rFM/QLxjtP0UDhoR9M6oBwjc3FPKfaX/g2aQNOuXsD
mvucIWKyyArkNm2Vpakn6+Mb0Aoif1M4vOpc2cHJWIKuCgiJCMciJPkIexNqGin6MAuZ5hvNIPOD
i+R7Pk0EL6uqn7bGle9u8M06BRr8hkuPN7lhB+4T/tBB+LvtOiCEgEZXnw4YZLXIu7d13m8WhcCT
NHlNMJl9yL/VXJgAXrI/kCut0XJFi6217SiYwB0BQEDU3/dEJGXSlsxVp4gfLq2fqbBt4h9oGFkn
nV8jGpUooYo4LrTqzyAPRll2/AwgYdoWnX2+PDmSemPxjocuS6wKADZ2sKhHDXme6CI6pZIjyG7/
7dSoJd5H3Cx03R8xODEgAbABNa16ZMVrkpkUWiXiDy4mtqkzlmUpXKlp+svTlwkOpHd2a6s79/rq
HajlQIKQxJ4xZVJuFetJcyouaXS/6s4Rm/ZBC7mIOamIg3ttOPUmt0LRYkK3c4A1mqp5qfKXzjRC
EWvBtvV5sxTtzhMqExrNvUAd+VaylsgtQnSV0D9TVjLkq4pLCf4WbM6hffvppICWLZw7osNPwiKd
H6VsJXx5ezicOzDQYfGu/bV6hdGosbaYgD7pR1lk7WwZZLtoweN0zK1LFwJe/MHZrGoqLr71r/MT
QYLzmy65CKQ2UzmGtcSxvCdl+ccZSmBlr80Dsq/NDxbaIiop8QFjTztQNBscup0KQuHKuYkJmx4j
yrjwyWbHSf9zDhtEC3PzeYw0vwYvEeqtV302O/dO5CfiQIvr/+0zKS5QJTstwDk5SerBor8SBRJX
ImllMlYjYk21yycMud6KReGNoSzQj8Ai9P1fnpzoNNHpAVjlo3PMKWDX0XoL9Q1f6OhfVnGBv0EZ
4NYFy/Miyal98i9S3ZAPYYDqJ0FJ/y1x3u9W/f9QdjvCTstX5WovnPN/6DM5qkq43Fhy7AslgCN4
A4ARq1vwPjFHb9CZEjBa5ZlVsScGFBdhhFosS4jOzip32lUnZ+uQYcCmUsSQ7wNKmAKIPvEZIoUY
dRZJCQN5m+k7oHZ1urSzuHNBODuWlFFqGaQQ4Bp5VyT+8H3XAYnV8BoXBsnZxw+0+IE7G9hpq1OC
gNgMTs7l6Hxg/+TlfQJEVWnq//j2jxm8tJH8MkNy326J0YhP3SOKhs8WG6cH7z+MOVDQWjQlYHZs
vQ+PaqL/hDC8VjvHYHU3dPi8j7Z33lJSrQXbxO3zThQmPItX3zpgGlHHMi1MDJJPOvm8i/UcylVl
NLKchFzZcxT+gzWWEfJUArBETeB82EbtHGvKgwsa/WmWPI23EQK2/49gPssH9DGPWvsb9fIq/6cE
RckkbLC8nDLFvkfm/sx3awCQykDONgF+txia4+GA7mB80qSj/rYK2yQc+EF+2T7LTBzLO7Kl/JGz
8SWHIenAQOLz8P6tdC/b/FG3tBBC/erps/tqjlZQhbefIRj9fhKji/j9SH7snbGCKztGIh2CGtJI
0w6q50ErAUxr0I5vzShJipn6AAmrHhV7kpkppZBZhM9CAyjffzVw9D5N5T7rtlgz0DGJCc54nxu3
NGvAVIlXPNa/Kc6T3VUopyyRmuIYUHDGex5P1JWCnaIkxn2OT0msrVFOR2ECYVh/ZsiUYk5HczDI
Rd69/KalNWNd7FFDpJ9c0Qfeb6z+zvZrHTOzWfS8hHm0yyOI4CnKSDeUExNua1ozw40HVv79ndq6
f26nQZkSCE1rOcK4KzMLd9m2YpWwtYaOgoEEUqr+qYBrxbxLvm28C45kytVSaC7FKRasNbNlxlMN
pXUnAAGB9kpWPAT/RrnQ0kCE7a8Qh+hlfe2TG208nx/9Nz//CoRon0uP6LtynGK5QUV285fjqo/T
QMe572sO6MLi3F/NzHTo2qTo4U3ORdkyQzz2RlPm5e3cz1g0jWYaLDSjB8ndNroPbcb0sfpTjKxw
LVpliAgLcM6tIzCx+eEnj9U4YmqyvJBJiQSOlvOqZtQsXWDB3S1sRHn1wV/E+edGMXoFeTJx/9hn
wRCBD9o8b0mzdF+IhAS7CN/ljE3uKKRHq0xul+ynsuHv586/HA1Ksg3zIcOM0fDIvcI1nkqFNAnT
ttTVJPOeZu2jCUk/4+Z/Mp/4whZUZMklfjKW/FJcW9X+1e5YpaPqbpMCS3EnfxwunZHhJ94cjyiF
bz3hkgxw9OxrIP1rHzjHSmLDSQ87HlmQwgkA8AsA932sE4yiu1JGfijhTNpy18f18UGuz2IEB3jf
Ii7E20r7DaJEvEyaX8f2q0wrGo3P3nD/vRkdANg4bjl/mD65j165aq7Ru04+40codLERwm7yx42h
XSHmaEiLM/shsg2RFkL24wVtsczH055ep7+9UZ4xjtt+cOrIG3vBtjwIvqMSdcoqowlQhi498Vfg
ku1NnixsVjmRujSpbYcNWqIv1JZQ3Kfoqc+wLo+BBBljpvEb6vCaIjiknYY7Wj33Va+Djidhn0Ia
u3Ws7TWowlXNvORBIfX5uyfF34HZKIJP1wQCjYSGv7YSmUsNeG+aTT8Ty5uPApnYF8M0B1qVneCY
AfiX8CKLBfimtQ9ILBD+YkWALBNEmmDkwphRr8JfVkQkNYOZGFhgoku8WafTcd5UIJEr59NlA6ay
QngQj6672RDEd43aHq7L1HYcTqRXVEwfwc7H1Q0MrtXrr+b4DuKdxSl3nMcvVJltXlkmXUAgX8tS
AgfP53lS0w19PQyU9u1d4WR9TZox9O6o7JRwEL2bslXq4SsM6bG/Xo0ShodOC0Qok/8YFRC/5bgl
zmRQMgCWHlBKfvZDVzzx3/9IT1OqxFzjGcfVMt9AxW2ttwppMWinltnEm4obWzRnTYbmcCh8SUoT
m9vaovu0tN2bJPTa6fNsln1kbb7bUbbDdBuKaoozx/bvXwYIGZEl7W8J9Ex6oqzASYNZrFD5jyVK
Quyxhx32VU5IHdfqB4B+RvF44ciHVZ+ozWZcm61IaXWPmAIXxy8y67P3EndTsfrlVrBRl5vC2xrK
hwLk21fP2qCEJr9pTVP7q4RRog7iHmiE6h2Hd86lP3WDIbf/fXRsUkrOPZfkv+45Qotqx/TPhhSu
60fQPlM6ibCowfqPCWuW+UIDDsXz6TNreGvrgmxUrqCHLHTKoQ6wHECqkXPSY+W/GrjrZIvszlWi
m0AkXGcA2AuZ6uaavqEIwkiA1DsPvjRGW54LcHgh39st7T/7j/xRyqNcwlsxkfBm3wfF2bc+wcmM
ZskxGAotVKX6i121kUFHpq1Fvd9kuZQqSWMLISZZGU+HbaH8znNooaLaFwX+emNqG0TKoZWEmVBu
mGHA6ATlERhN7rY8mF+v/RUIJgK33ur5n5/+rQS+B4h1azkq54bQSszJwwhILg6iYf8+MyiZUsi1
vutWox9gX/oKp1ZlS3q5nO+NXvl9CxjV9fwTi/neGQS3jvlvuAuL+/fZNftdUJHx6X6YnrtnpMZ+
B6d6U7eeuWe+PeTUCQvFmlt8bhM9DnbzqewxynIVJesY7Uov9GGTbjk0pPS9C9FO0M6dw+qSdrv1
ZUDOPu69UXGxNZGfIX9QBBWr2HNxvzpgtV+h5Y8h9Fxa7iA5c2ma76+UeyC4zkKQh7G+UU3GiHTb
cJPggyGlC32i0ul7iV+wRzP7FwmOfcoxaXT3X+TgDm/TTjWBYg2i5AhM43CwskwpqtCfGxYpgpj6
5hk10EveEo8OEWWUvzsLbZg9iH43J8FyUWK0fYgXoyFcBT3uHH6pTkk6+NeJEXbYyFv+TjZchkUl
Q7E3k4nMGHq/ERbESAU+nUrbgohq+L9ueqjg4p/bfhAQVssP18CqgPuICBoV/l2hJl9Ub0P1ANz9
2RdWGQD0LdiVt0iYkqWcOzPn9lXd8Ee9UrF8xbWX0v//+OoeSVjSqeS8SB9BrPiqaHxWdFop00AT
P8mXkRXZz9LHM1Uo8xznN8+IFsp0sXdfuaoUYco2GXB/XwYRfRVyORWilj00IpHLCmXz2f+sKtAV
evaBC6C56XhmMuvAQC04OsB9STw+CSjPVfsN4UrYMfTJQ9snlxpokbL1LejBKb/L+/xY3FMTUiP6
qAp2RIQ2K/JbwVJmiza34agWwpQGCxuy/yLjEmLu5NdkIUqX1X9v1hLjt6LQr+bBMd3nSmpiRlEZ
jS18kdLZFmay8/2ZZfe3CAfjmnEcrC4vbW0yRD8l/cGWiu2wMZPUGfO7sEKdZzk1/kpOMgiUKUhx
sHaQ8JKpsT3QUbP1HWBpR6+nwP7z13dS6fd/IGGJoDudbadfPb6kVoyj6LoUhtHKSEn0JIedgKxr
urQWx7+fFixw96ZhIukVtLKPnYmBun6OgbUPjfiQyCoAFBA9X6p3QM+ACYBRK/cqtL1BpB/Q81qv
6MuFffbZ7i+VaLWMqsVD1yAHuNiSvYW5UwtKEhMlXDYU2i7l3bMTyL30TzsV+/cn1k8BTVE+hKx4
s9OfSNtdBwER39UvTZZMl+z8QKm3KpJVHCByTTIFzSKds7TCVocSvLhGP4HEnphxqOVe+rHaqGmY
DdCu76/zA7TNBShbKUvNg5ONc0/DHW5EgWmBo3jqsw8auEvWUXruXl/Xi8VQg6Vw3UUFfD5ztMuk
SfHxolOWqrI86oMTineX7WGZ+Q8f+izYjV2/9/qdgK+a+kpJ0+JXpf3Q3AaqyU/w3I/LR6B8Stjj
HWwSAO/dCmvi0SdA/b4VsrNj5DYTcKlMsOzqBsH1kqNvNAoFU+O4nUjGVSQe9KNqRgvYbMwfkcSi
CtJPsenwFlxbN2Y9E4KRXD/1rZXnF2e0LjwO8wCwFFsgl12GRkgjzTX8J7Y8aMmQHVVA6ZBgvq4H
Bdjii94QfDTaenWmRP95KM8cBkqCgUFWa38EwyLauL2fjNpw3CBuzTcPDUHQYv/U+gUWjRnLgqQD
SwZz90u6KeehUSqLKve0g8idiyOkAdnPFoRvFOQg3KH/O+5S4nneHV4Q9eTi8Ta/r9Tl52w1w5rC
EmIvpOH3JKRkTHP9euhQ4WfW7/vBaXrx/P9jPTd9lYfZVD9SCDosKr8nPNx9aao4ucZrHUA3Smjh
1974sto+bd7Wzi75i8EeCsce+wIEf6QVLnFwtgYyQ2agOryNEs3xzAO8OPx/Avcz3qR0jqS7a7CF
C7tkBrUwt7nPOG+Yxcu5ZrK4XTg3NwnE3zRr7su1X01g6L9eMUbuOav+7Ws6FiQgz0RHpVkRK4+z
SVXhVmjm30xfalvlvDjc5B3YtajyEaC08C4Hyx1+MFJCPMHKAOSZSHcTdgw7+SdriGByP2hSSsiy
4SoVMTEeehL2+U1EQzAuHOITL1Rayc9zKWJJocykN6U8xCRPx086B40pI1CFhe5jjPOrTM+GqV9P
tIW7AAHIwP3nHeCYbTfYPf/LTVA9iDw0hd/3boMERy6QB3PaMiUcWcJOi7gCQJ2cxOEUgZ2TNMFE
hO49Cqosed+++8pSFVN5oVny+mHkvRbHrhdw3L0tB2r/sAXea6sgaI7+Cqqiyhr7t6SgOTJoI8xQ
PPbEpQsypbjUyYVPCEwurdAT7AFw4ekqecM03ArsSgfacwjadf8jw7nqVUIP4MfwM/oFCpCPwjri
oJwXKaHWpootBuP+en1sZW8xNhkd+ROy9H1NB5JpDdnJJ4FQoYxZdqVZXRzcYDpfdPdYL+N6ciB+
u3XkKbxAkLtuxptFXRgUBwaEeQbXk9xmDaMkU7pxAXHX8TVvu5YiCRhcIQ1PxQqmBO31rxF1A6oY
rLQkrjBtPJ1AqzOkhLAIvkCHGAlXeb99+5kJK4m+VD1aUw++q71P9KwbkH4pF05nBuYQA0B8DcGW
tmIU3G2YCyREmv15DrKS7luEUw8bwyxnpR7H5jaYPy6XFUvKjsE1srAIbt2bC2dEdWpLl7OWOvg0
FtUWz9AqIrD8SdWpeUoDPs7pVrDL3GPdYuOs1T/1v7zuyvudwkJ11YTdIC4FrmlFz82eb/Vfpf5x
FbMmO9EaljrY2bnSkiMIe2ykrGQh/0BQLyQgvr2b7qoe5FP7wX8EUrTYhHRk7IZM2HOrrmJPhtwx
mM4gZwrs4pgrSuz5ai+Z2AMcPP8MITYEaof2UtytTIWqgEZQdLKJ6DtfJPYOOIpfExsU7P9wHCIr
LpjafoQPCCsOa5LD34ZZfyuiuqO43wS/oRt7HvkHnCPgThrsE9warxyEtwY02HK3FFcyTUwSalak
weRCHfsLjLB/fHQfPFhtt/pSoHDNnqcEJY1HFTStnFnWTJ2FsCnoe+wpcuqX2PboK2liUw/nFse6
XuMsWZdPIP48VYq9KApLsTrw6SycP+8i09K88GgcIyW5BMcks900GbM2UTbhSsbIRdKwh9YrjhqX
mk+YnVi1qSQjBlVNn5r1ODwRC31LJjTPiRfejlhsn/M1+drtUXvXmoNliS0HSix5ZBObbabZyL1T
5abuEVs+t5PPcZrYGyBp3royRaH5Q90HiyXx1UIP3cXlfT7xEb9b2m5XutQlsQNbuJUw8mtOYaMY
l5ZYD2Mwtpzg2TWAyEo0njOnuJafX1k1zON+qu8YNRNNf2bMzV2HSguKzRuOQ2mz+EI4l0Z2lFdc
bN4y/dlsPNSs954amUb142LIY8PxMGzCImfaz4fdQQ9AVUFJGaSkSpfAZosTUVbBast0vxyBHFNZ
jAanUaK8py5ZVTeUe/o5VBEiRexSfHWe0TC887nEyjg7vqZ8LMZpOJQo6Y1pEWxxqWrVY8gHpm0O
uxcolICnfkjc3tUKpwYgur/edk2oH8WP5235PyC1AyLjttQze2oaHtQnPgccd+FwRhf3BAb6VlE4
ozb6JUG1rzlbfBNSb/DdW8XHtoErTx5z8RANs0M7zy25enW2f69r/4RPaI9zRWbtnr0H5qCl/eWT
XGpUUO914k0BL8boI3QDRKpRR7WOEYv90LVg4nbgg+4PqNtvs/zW50l9+66kDQUM3pKDqvVwZ1a1
6O/7xYM5+Jyr5atEODXa6YHqvZvUC1SOSQ50eX3RAFq2lZa5wbwrVkgUkYGHqnLUeBjSQ+HhKe/S
CjSi7m0jSp1OySr4iZ7ijeeHhGUEQHUnYpJDHICYkfjr6kfRR/WT+rH2vOIh9O6x+az5AAKQiL7P
mPQHZWJIoguacrhX+vK7kpXt/1sQv3Rui9oqVb1n11CXjpgE0YJDxy0NOcI+I1AGO9tJ3A7amcY+
6wS8sZHWGX3E5m8qLX5mmo7gURRv6HtRas56GHtkL+apml50jAPUFrSS7RVSi5/urjiMlb+C+qqi
GslmwH0sKBrpFvdbtFFzbJe1b8N3o3GCzyHC7G8tkZKO9QPZu2jrUupz5+xpQ+W8fLJEzL0v4c8Q
e+y0Ys0UUezcIPF+E1jXUMSyTRCfL+znr289quLEVjwx3D23ddJjiTa+0lTD0Ev9BcJwg4xx8u2u
sxdX8ZxRwDoGl7eZ0MDU8gmXY3WEDtJC9Hil0lCY/4Hqvd+TE8/cXoqFV35j5PE9FNXr5HBMWO8D
/BTm8tkiQVjP6LCn2QQPrTz9FYVVdrHhIYKuf7XFqwn1KYpP5kS9gJL6i2dR2o5SglW6H43JAwYv
2zaU2vCr8stPwRaOE46QERrWwPXw+WhfHiVy0rh/gtH5sfOvZubpAdsjnAltsMeaLf+Uetg+05Kt
ebWKpe6pEELiWHWOR721+t9k3T9c2Sqqv+drnr7jZkIR9hODM6Wn1uTS1hNngW2DFsav986xUj04
5fRGKwJuJnSNN22LXqqv+UDknj5ojvOE0suD8G7LDOwRE4Gl/EBJZlNFqVATOtflZxEEMdqHl7zl
df9y60TDJYCVxYTWUUY/tpLxRpOA9Dj7J0asz7dsQMUKXKyYn/KA/iwPvN5QV6oe3BlyqNbhdqwB
VHRknGYr2VULT4rpcUEDav/BkyGTO3NgpPxrIQBRGhsUylbvegGGzZgSmCb6wAVS6PzyytOeflAp
oJnBPPothQx3H3TM51EcZbxOxduA5wJ1dlC776BlUx6Ib+IkMdO29VmocyPK25n/QDZhGAmVTkg5
KjXeXskareuatK1OhypsrSItkU9wFFkv40BVaV3NLPmAO/VKiuDDzhjDMNRm8LBzDgqWWbtT2uC9
ffNzfE2A1uuBDuI0lUZUh6PPmxtDpUC6yUDgiRvgbqiLuDojmzC8oE7U80xadq3Ef4AVjFa7yrYa
WJ9qlWI7Z1QhleySIUSsXBZAbI1Tc9JBmiNmGslv7nZb2EfwbekReLTeoJx5pLGCQcEPrURpv9rd
08mqGz4aWYIrKtib3BxF0vkA4uQ37QFGyoKjIag3YmYw83FQiYCscavugCW1S7ctdXm06ouFWxCb
0RpzHqY=
`pragma protect end_protected
