-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NuxCXV2RfrbI5cPFk26wv0dKXvbAdCel6JIiNmoLAp43nZ48oZsAkkoIP1Q2rITGikbJxLc4/Gsc
bczipMaK9Xr6lZy3MRta9Xp1+kxuvq+pwamqHP/R9fekEK+xCxfipbsbVDzEIhpRG1uxmg7MsltJ
1FAzpA53qydUfU8LVnU5DrvoXMp2nsWIJVLYiZ03xkMG6860FPOkbOXUxhWXpXOM+o26RWx8cKhB
EZuyxXIXBL3kxLbEMsfXgJUzop+P2GbeRmjA75d8aVb2kDyIGfIxnIBh7kqQK2+q8hzTdP6YTyn6
WiKPTLiQ96kKNhRURZVMkhcZgLkmY0cAcEZDQg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3328)
`protect data_block
fex92h6d5MSUq4t2uaTvQ1xiOMSEovWAoLyip0jbVapKX+pmvrlsPvoz+zdTnH76SEiLcEw9kPic
ERqBH6DOckC1JTEI2u6PybyiSAnGVoeq11AEi3AIbvlToEA9oPn6dE4gTFZAmRgydJQwEJqCipcH
vahajjGP+bM/oj+2T/Y3Bwq65XbR6WC8H3vyFpTbrwU/w/4Qrsdj8Oa29OCA9JWMZ/ixU91ONJpq
GpO1C5Vhgr1dcUaEjBNTgfs4cgkSCsq3QHG8nmxCtdZHi3mIPqhqMJ4JJlHNTZNA3qyJVH9O+/sX
2WchXE6IKwsSy79B0nwdgX4o5JKiCrz+F+zp3wVEGjzKkxgm4VcehOkoFr6YoumsMpOrz5OrWjT5
xngxV8VMN2J1P03wfHJVw2G8Q0qaqlB8pNY/9AMJquQlo8BOo9/fYs7zjzI+Xbfjreber8QvUbuJ
SAgjX/T/n3bP+2UFqLAVKEnUwqHd8D21iC+ojxPJtr9BWtrbKIISrYEUuxT2lM40b8RuN5a4Nu2v
lD3KXpm1/vtOSYigEaB+n5VCHsTez9D3QG+zCo3XGWpvMhJB7IPkYevbxd68zznoEcHk5L59+J52
YBaCA64f2OxQsWbIFHN80iBgvddWMgLTH2LfEzGAQRoqxu3Gg2H/DxihpVRXUqrDaSQYp6D7xZzD
G9oPEG08iIp6/B8u8695YFKHHsXa5ExbfZCiHV2+Yt66mObdboHpO+bKEUy0zv5v4YHbpA5yfGRq
lM5zZRjVodiLrWIeHBkyRO5M1PKX6BrjIuyyrO4GtstiX7vIMGWlA5JyJlcJ1udbOo8aqaRSrEoX
p7S1TqacOtXg0G74Cfyg3xerYf/RPLnNwLvgolDMEYohGX0WOX8Zli2Bpr5aEmZjD5fljUsJWHKL
At7q1B1KZI+snhG9Kn8ivdImafI0G8Stnd30bag62OuI54JO+ecu7FpcWZEw2TMJUr9od3t3qBB9
V6CN4WYkyAZ277RXteaV6VZCpCdwfHcRq9kgJDosGs/+KElxNjO641Z/O3X6F0WgJt0XWN1w0hZ5
grXTRiiSDdPZlkFd7oEzPt5lLIhWy26q+wd2qK6mnXDFzplXP/zVMCSdpouKzNH8FVkXsVsLTHlF
eKz3kMSl5lf338tErtbmhYlKv2IVblhrAcZE7rZKrHb8/ynqmqy2qFvrR9kRx2HFaivY4Nzrp8xQ
a7mMmJ9fO6Xicg1s29J0vDEdfQNvCZTCbXT+rDJu5pwekH7Xc1T88dw0dqH0L84Am9n94nRWJKQK
CZqpQsgTOIMEhnzdWIzK21CtCAYBQrKidRPcN7G/SnThveoobywqKee84k+lqkgEvFaasVX3rv0V
LgY4ps1uLrueYQCLkH/474n/UW5K1ubsBjJJcALJhPX3N2BUHnhLdHqZWF/8+lNyovo0c8Tt0iLU
VK2KSPcjq+wl5+/CJ/Z5dWGbGGsgi0Y2YE4etld7dfEwZxRZgYTbocyrMZAAdbXUFXvlvZknQCRs
VGtGFK179HA5jjTKdcSgY6Xqwl0MXFI67b0Rkd9EPDfmQGnvhzrC7KRwkSEcjkYMp1Xb+rD4/nJF
W42wWhbVvqWte2KIvU+DigEX+qD/cjwSveQ3dNV0F1a4kCs/m47CMRHkIRMZg1SjfNxOGgJDJ8cK
QOb3OEEOMMH/+BrZjhoe5MtpZ3eAy9UHxxq0eYIOVx4tknZksPzGKNR0CtY7rxRWCgTaXZ96mcGA
vZQpIHxJiZkSqqf5ecADzbYHUUqfiJCoYvAWYCt69U9HU2bwjFVUYsczMi1PkLIVXACCi5cvhJLW
Kh7ftq3A+XVxQqrgFf+hgC3ved0BmCpT7bmUzLqPBGWEs4ulXSX3N8lNpRef+2C+MwQA87S//aaD
YK1b0KmXTS0vdlyKt99xpI2IxHLDTkQP4Dd0ber4wzIwsldqvUexUOidbY4IvqGKRZYbLycO7Jbi
nlG7I8JjCY4Ab7MfyZFkGOqyyUCfwXHW9vRsuaeTnf0aR83Rzw0agrmdrR5sVx+Gj9exWkcBo7RO
2+69UFFc2loVvIxoBNOLDM9uvoh3wwEwvH5uYwhYy45f3TsgKokS2TSXaHlZrw7hdnH7qLdwa++o
zt6SwAlNY9XcOjwE+v0CmvGcNNsP7dAKD9KIzOssqnTNQQXEb0aGz2yfHV/idmVYNnUaS+fgLVst
zF3v35kb98lDQ27lS2fzmUgrLgHk7ySgxXtT8EXppSohSWkmEgsSBB1XMP2/wKTSQUG7PpRzQo1K
BPL54AsS1RFq20NxZMBTL1kds2NOizeFM/L8RMOY32QDBKDyf38+b4LUiBwqmK5v2XBqJcC1yIiw
VwyV+B+ltPTRg4baM1OSW780tDNndk1Y5+TOTpoCm0QKnzC3n/nvkuBVKMcUcOB49BsTXlcBb2JT
Xl2SS8v8TQva7/DjjXfuS2f2sIe9pgYm9H5EnUj/1a8dZquCllUyiQJcBAZKOFBoTt68EbMddaYY
LDqnCfFQeYVAMR5VAB1tENwKfakk9RW9WXVUc1G0TsTzdssV/TxvQ0Cwjmt22IjuCFmYwfNAapev
7bYmoFUlmAiMYHKwmLKE600iYL6dyXsB2J+xbMxdx6vXAPYxKI8HtVXjXcwIUHQ5+QGDejZh9zXs
Dab5OewUENTaWsRPr0dEUwmXjqgsJiCD2Ilni3GkXyViC9OZlAbPyTw0PBWsILPot+NAlIIPGjTa
jD4QrrwqaGsdKoWQ7DEUqJqGRiUQWQy62J/706rA4Sus7e2fzOrF/6T4rwci9t5ZsYXMNjre+cx5
j73l8ooHpI4osv8PiLdiIUoFB3Gi5I93PxoWsQ0g85FCevU5VxkLOkMRxc9BQUTVs80ZFmIYF8lV
arIJhGve2k5/LlOjqbSchT9yWplaD7gB0bnJZYKYLdGjOxA7ufFpJ/UO6ELUqSf1OKWsNkeXJxht
5JfupIfQm9Nkk2QHTryUDTNEXQwmQPRs9FoDbavS/zPHVcnBGA9B9KFNveXYvLM/5A+CkYzN34Ua
3AHswKR0glS3eULlm1ToYz2lW5KZ/lgVpN4PFLOVIrRvVDjrtD46qnngL0Nb6Z+hHDSDvbScYJoE
9p4hA5vB/ImhyJloCxYTr8UUzD1f0bCAtWSugaymcimdXoshCSUtR9sdSktIDkQTDy1cokotsAdN
9B6WBxDfN1tKkLpXmyiqmgX+w+5mk+VTr1WMwKxA8TGOIRSaD6wnwmoFa71QirvsFxoY5Eg524uP
GAM6Oi7aOQKrGBCdMNPMBdPAC6zmI1HUcFWuX+93ojtAzozFOGWo828JqXdb4RMLltBzhng3JTPc
DXBuj/udEbVzX3LApHVF4SORv+DHicEvVKEicV2al1JPTDbbQ1Q+OTnCUutOmMIOqpuJdUo39VLN
viHnSw4y0h1FdNmZjYv4ArmYRaG8mDTyqnNOpLByebLkF0ytxs7t7f7V8Xbx3nO8euIsP45LEdS+
ospJWgP3CJlrVDrp/UmnZQBiWVxBWqaefDRzE732UXAc2h2zPwqXIzpDqKoi/v0zdGbEA26bIudq
RLD+X8jzNYgRqoWA3+yREez7UBiye3WQifejBE9yEsXGvK8troTVd2EGdDRpnbVI0vyFLwN1fj/+
PoWHeO2nYqQ2muF5Db9rxppe3/rzcWCiEe3KjtBAzome+DBOQ4edVdS8PQLFFmpGgwdaEzP3gD8m
hemDmFYVxHqbzRxuqBzZnsvRuNrqdyDXyqfUV+suV+62HtTU4lswtRH2JUId438y9hCw6cPT/3on
a1DQh+wl9NgVG/mrIJpZ94M+AjPDDLYXuXy3692PA9k4R8veYS51exm1Xem9O40ncNv1zUAnglPa
a2H7+cr6JuwPw4Yk4b/OuI0jnzHH7wm+gHuaC8x3g4TijdaloYcSmpfUPaWA/Pp8HIC+iI9YSw3W
OU4+DwVWtPnQX2y9U5hAs9JqQYrFBZroGNlH83maXn53kU7qmbc23dNrZ/AgwZDTP3tkl6cl9r/D
Wxpg2mx8FjMaIBntMBwuenmMtueMpK1hUG3gEQA3LUbnC5RPXI/HGwTqYef3WnhgYjoUsI6qs2FQ
LxsRQzJtxwQcqN6snXZlhIOGQAKp9P+7lG8o/poSBUF0CzM+fdpQOiyxXGin55C85OtC3mnNNAfS
eHVJvGbUZxObY3hVXbuLH9utwj4+BDwLEGGEbMoPvOIHSzrpE7Zautoq35EOtmMbnCzJ6jdwU97v
n/Du/YmnVBADvgfHHmLd3kDqTH17fpIAK0UB6xa7L2ywid1f7MG8HejXI5jfHkiUnzrd5YfhuYYX
/gw/hdvzYKKk3NLVa7W7ufYtV9zVTzrdq9QKgYr4yGgThMsGlWJtV5omzZwOoyqodAi9fCLQflMs
D4Ego+Clwn2EATXFYdFy3v97Nm2kqw==
`protect end_protected
