-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0hqrxSN7/TjYzCfoIyajTPQXFIguoyy4x0mMFxi8bPku6nv4s7Cj0OCkfAyijb8HYGFmzbyZUsqm
/E45KCW4pDOSPhls+dcVKvx+7Ruo9kMSuNBEYsHIgge2uvrBzv7+ZIRwT/T/moH2ipPLUg8pSObH
HrH5dxNQ+Ouluu5ybscxVUcKBQzScnB0gtfLQEC1SlzV9nXDx5IybpK9fefXS6t08dvn7rcLS8Lb
I+rXvHHfWYtLzmZ1FGHSm7UlvYQ5TbnErH4rBKKESnMyigfj2uFZfro+phoGtcqZTOcSOcODd2SS
BJeicRvg6RcjZJjT6k9/1KLxXDjZTlymW8KRtw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4528)
`protect data_block
kbefFG2kCAHvxtkBWTaHP/cpbomxfgjH7dTh0glHtshSru8I+HCAwV95r79Iuw8o0HzlDWC4l222
D0Mfp0Xoj6axFYRbo7uTWYbiKT1046GU2fdHkDJXngOCllgJDzr305oVnCkjYXOQjmI3yZlv5R06
zlJ6dqOhTKRm5tIDtNiKcb7aJL4nqV/fkLvilltl56r78yFJLjUWdlOfrssnDRTs+H1LAOYFBI7R
jxCvn/H7X3XMYOmPZdnNjMWRsEpyj1kpPXzkuYYeJPPzuoM4H1S5uktkTGcyrazFnX/4p6FehW8K
ZeZZXBWCc1nahCbNt5i47GL5y0ItQ4ekDRtHkhITSXsSQdxlofSa6WLx3VXk44XPK3cE+sS9+1Ii
EzkYI0rbLd7lP8u7udap4SMYJ8E60vt3vsC0reQ2g0yqCXZ2TdsNLbJ3KQRpflqayS+i+Uit8vO2
H2k9/8qXXP0Wj8LJ+54952GprpPYyfuT4J0tt3Ovk+0Rz8fa0+XJP+mkNSdVjuWOEqSKk3EPywRV
7BApFi7m2ADdGTJzYnyzhGcgI92xuDMTO3zs3xt179+bWB21A1YxqyTgpiJF+neN2PtCZt4nb7nh
vmpvsTuUdpNfUzqRP3GS3btZccaz8RN+ptLRsPD2EEQMXcFrrO08Z3Z8LzadVN0QjGdvAdlZxYQw
R2RHWOYNNRbCxABE+vi2BI309tBsnBwW7Icl4Z1+KiQeIATHVha+DeMUxdYb8ueeUQXRzrmQvNaP
ctJ+wfZUH2jKVbUCRqkzUvPJIwTHEtsTxlA7WBeM8grGXrByr1v8gyR+sxSGmwojHTWqlblcx4j6
rMkQvYf3Y0RhJ5AeOEEvu3kj6SGkM4tdk8l4ET4WHVNJEWYHlGM9X0amtycou8WIvl2ryVdo6wJb
GEE0G+M+ff1sMh1QYv8MaP38qk1YrzHyUcEpxb8RgcBz6CPSSRgMasOb7+kOg3uRmywXpjYEvQyL
v5ZhdcykV0wRzg5XvHnzP9NytY8f8Yi8sz/k8xEcFIY682l93wOsB7nNIM9rnYS+stHewD1g7Y4F
NBXY41S347y4qP4yno627+b3JhQTy0jENhrU+FfTf3j+xmVcjIL0+X88Wd1Woz/Lqla+nOyhPJ6C
teTqUqR/xkWCf2LPxlVwKxVd/72gvDfqXrAs79YKbrnCYLWoYT3XjDusCGGAmq3f/SvLH1cgW2jn
7Llaw7zNosL0Kb/6zWdt4gJ+0Udl9HR60rRcXRti20lRcTiLtvmUViUY9NrgJcQH6GpDYY+nsBED
ux1bVMbfmrBwCfzXw3b1SYTB4I8PcY0FQ+s75YvjJwAuJ4WJok8T15tHvkK5czeVuC1jbBiEHmNK
Tg9txPskb/ZAftJR/XLlaN3IHmGvpnKW49eV8nwwX7GK/ECXIrTk44N4L/LlQ8DKx2j+ngAxJ7fs
aKL9sxTvTSUwobTxY3KSUO8I7/hY1eObistHocnmwHN+1sNVd45bYOsf5hzQn9onNPQyXZRZO+kD
SZhnkb2CEIRkrgR8TuFcwGj9j1hSL1UxnDC521h/XjZqv34cttHipEXSqd8XbotDR5gmq50TOZPu
OpfPJIrECDt6RzWj/R/OMgS8owNXCzVKG5XeTmuq0KKH3VUHyKotWtzmucuTzNEBxCpsivWTzNMo
4RBSLfGsPfplwGQegjHUOSCotAiLU68vNN+ujs+1/aeHBL0huF/+wMqAx59j34GhMplT53fgCLQp
A88kCZbJ+MKdyoRs7gJ/0a2/GrNVKyHIJLwr/vJnhQyUFe1qje/ROQfpyjNGzCGmpZbc2Z/rAd1h
Yi4y2F0Y0LmR/D5G/Te8i/G0/KauYijbTvq0k4MJyuJWv9yT1Y9CKSFL1SoLXJjIUzP6IA6z8Skr
Kfs+pkDN1hAnF9Ghdeb9cFUFDxivvvNpGwWe1Vw8e7VACZXLtQMN3aVA4nsgkzHGsDzraewOmxz2
6g7voV56FqnyXZWUf/2fnJNTfew+O/uNcpz4XkJf3+dCnU+tJXShclz4RelhdTE1E6aKo/7Y2TtV
YeR6MzOKEXcYToBran814QdrDVbsnFbgj2PFjEkoVeFvdLsJJeQQF3hzthhcI61A2fLX8sSfSuLQ
SND/0RKjlcUUmVsSov1CDgxz5oUEim45QoDB3UjnZuXCG6mhmJVGI4JkwjRmaEgXO756ylOtL/5p
wJNMq+W+itkfD4x1CgPnjyT1yM4b+2Enibd000ATgKOjyIPJlnAZbEUIRF9XEAvJmQJmzBqvRTrn
4ePqZDaY3US9AeprsG7ND6dDA/3rrkWMmhTqmnuJiWeBqL6/bbgdjJZ4XEvKwG2rB2e3aI8gE1MT
c3YGPPbwsdW/lislBkP+jj7eMvsgl7Icd4X54zPWGbRP/8M2mwjgDSf1vBwPXfJNQzwxFAxTv8De
5owPHHT8y1pYbaPe4wTtEaaPfz7eBNJmsXe61Jb2vQHZNmSI3sgicvNmQSWbuyNWgx0q0I4O8Unx
beWPlaicLdA9WtsNl59nVTLqCEXYLqtLSn2IiC2yRUiUDVRH/OVrt6UAmWVEuEyrPkWmNYw29rOF
qf3ws83RbOXVmzualx8B4aRd+9+vu0TxCWG6DBH9/1dtH8zCWAd2I/qaFzuZBFYTATBt7/F5TFDp
ydyVYs62aE/UMl/LDPQVDVjn2Rh9kEQBNwQjpU7MihACU5THeJTUlrKS25uJ0cVHEymDZBaYpPed
kD0mF//u36PBDvrpaUSMXugGalK3K0M/02GNZzstpjyclajYRhX5RsuDi+IP8qJZ3fM/s8NBbFCL
k3apNXdlXOBMrG9FE2sWf4qc2Rl54Otf4MafA0lT2PFvfjsY5I9cIlzCzPqFB/P5gQ0lb+aIxUQS
G17EuV8uAzEbRLyr4+PKlCrga9tKkRUHz3TudxzW9Ot0+RIw2cBUlgxUoaWEhy1IvRvPe9of8g6a
vxmu4lt5AmTbZUobgdwg66aU3H3ct7V0qHNv1de6mTCPVVG5AfY0k1nIO19zvRFlcAZCz8a+sq43
esx9uAhwMrq6OOYCcG4adUaORYQYVYopE392BbggmWiMoRVlLVAbGyc1EDafr+TS95QmGU1KZ0UM
wBIr3vq0mD7h5NwWede3u79HJATuzEtYP9ybA0dRZj5i+hZYfrMjW4OLJ55d0QSIiwas34QM5wWb
rbmpALJh2nNAQjdPTm31YuMtI3xun2pO/1s9gk7ZDfo9m9E3TBiVLkExRlxHisE/3z2PVvl9+az6
71bz/36AG9Z6XQfTUjdru658D13YldPRwzbe623qOOEBgMI0n0ScUiU5Bpj8PdaZW8QeatKoiRwk
wpdJZsFadKJWV2dXOy8ZbYvFIJY1TW2x/IkX05q6qJc5zColvP6c5e8bh+nAYzOSU9glIy3reJwJ
z3bMHHO11nQfODFDy6OlgXLdYfc2WUpSGeYu48YFm/CNJ+PMPNF75f1iuAPV5NnD4s0dSUCjuoCh
o4CHpCZNhjPLtI92gT5dNEeT9/2eJXPfebP/BWtizQSlSc+AuaH7zQZUKC6bV8kDk4vCMoJxi42b
bjsH+cHysPdQ2+SXkpKGhlcdwPf0qOsmsq4uUcWN1mLTnGIct+TCnkR5TMK/uSFA6BHkhgCdPFFG
xIOK65o6+NLTCzQ2WZ8p/oFmqJcOhI8UK46K1dGwZZ2EtAwcAl+20+c1UVXmDtwhtycNiiXNwT5O
Hp2jUFHvr6F1e08Ox9VoHu8Q9+mITUF+LqclPrzlwOZt7F0bQCXO06nTcPjGT0E/2QrMirqqWcm/
jqqNQOSO0XO0+YgrbElyh0B2ByQOLUsyGgG+6C5FZTBrPRAv/bRTsBRxi4+gWxXXty+jb0HYFd7y
3J8e/wusuZPeS5BnI9H+Qs3mJO7rnLaO4k6UDybioNomQwtdNyEs/uB/gJO0tgfNcTWSzGhwl10G
DEs/Kzx1Z9gLzS9vj7KGaqxGfFK5UpNJpDyWQwjoz0irV5aZiGcrex/TcI+dQ+AUlQ0IQsCC1D4c
oZWJdxwb7T3f9AAFxiZpjnHSEfUR+9hzfE/bMasvCjh6B1efnNRlL6F1Q+ltThYtTHKUYgCoKfkK
2Czc62k71EmWg4KbIVheceLhpMLB51BZWVB5emdVvKAAHu6MHF1qeDkVZWVwW41jGQiMgrdKIrsD
yfsIYjP3g7g+JVYY0mtG14RdUZciVKJtqmsgHTHctDMdZChmvTjTTa6jZsYoC7MhLnu7e+1Y4Wi+
MtmGPdMuGq9b7Gp7dZu+Ho8wSfjV5cCC9Zqp6oAmt3bp14vOkktF+QzhCLMXKnBiil0oBywIE6/Z
6a2S5Q2io1kEj9DrCJLFagCWoNB5TMDm6ub3YZOdqRNUVHE9DgQobSZNQW5xV+eX6tUY0swaJSv5
QMr84lBeRrX8aRArU00/Pnmiq5n59UsRK1FCm3LTamUOjU31KKqvI1z/dj4N97UzpFumPEzbNWpe
/6pqb1H+FUgHv+XVXRp+glCGxY8oZF3dqluXMo1F4vH0l/gClLZQZQjTJOErUCn2RV/bEYy/SmSs
HcUtMi0+nOQI9hMvxzX3mQnoVQbiTHEAaln6y3o7Jz6MqYdCiQ3EflPfrn2kUc7PGOLd/D+VxUBr
+g/r7pczBQx1n8IGnq0mUgpwzS7OVn2pAlqeW6uCsuGHGPn7MNmSVZa5Fe0DLO+FaZJVN535hDhq
//iInNXdT1IwdxgYehcymUFG2Z5BO9ddIegZirqxtlaXpRoqM7tBWU3G3MgcZRNnNAVvhBwGE/En
lqUKNnyUkKo8vridgvVaJUzMscnPBFcwVVw+QcQnAyQwTGigt7Yt3Fo7WBYHzQWlh6rAJluw7vcJ
GcGM2LBiW48Iad27/RZE5r6hJOxIV/aOMyllxybpi5ViL/p1QtA2RNi+TyPvkyFiiWRJwKsn26Fm
INgZtdjWMP2sIMpspk/6z4yVnhO8mpH9CX+g+uHP9XF1JS3SMonae/Oul8O8SES5fDb2s0c9YBty
CpmtU8rACeaod2bj/CyUasVq6hL5W0Ll9MmGI+E66yWk89FIfrU/DHcXNtYZPfWMl8p5LTjVqYp/
SAIG/7SMxXkfpKjBJpnt9GPl4zsxYTN7JM7kK26nAdLreuVL8r6H+iO2BK8+uaUhSX21RFvNPMov
70VDML5eSmT40Rax1yydm8QnDyqtUBhOaBDNwQHDoQx++5jNT8E2Cb4VCsAJ75a0l7vO4AdRgfti
HAGfeK0wEIyaBafThToIGEcs7k3i7Qgdu49krY8x8L0p6RngkEuLKkniztpxpUJAvJjmpflyUU6N
AYo2aA2rBBQlThRP0Ve2ZueiUHN1f448YFlcvHNUt+gb92PtHirWFjkxeisdhFFMf1djIhGhcQKN
wySiAZbcDWTQV5k2xf1hAVLIJN9tPbcWzmG6wuRzjBPdlpqFG81KjnSqmRbcXBTEC59P2co7spBx
NJqiFcRuhR0w1YX5DJUMrbWCV4rg/VRlqWXc/qpsGh0bKArb1C4WVz7u/LBunbTMPhu48tzGZwKj
2E433RJs3Whj/YM70jsboePxut13vm81yqzqebgHMA3Kg/aLNfI2hxvz8XD8OfDenrI+ma0v+h2h
lcw+thjHhEPJWn/3Gt+HfG6A8060nJYLAGrw7mN+ZpHIs8RJGRrfqorCYhGYm7cNePWQvsLcp9nc
DIN6YkPKNDBKll0ojcjkjAELUGL6W8OW4ZpbqwweorIzcqzirkCkX4j4gQhpuWx/1bVG13B5Rwth
bkEYKlp250/hcmZSvTLy9oyxItniQiwMl4xfwsDubqz6kGbXlQR4ZMEW+5omKShVe3yJpByPu00G
8W0O8N5o9JuxlanBS5m8mzxBzZcPQ5Jee+8/JNrt493Ij9fRx8Fwnen4g22zybHhp7jrnkW8JQcK
7E9XDZnk998cgZ+tMVtbL1hwHf6JpqMWwfZPbsSJeohwg42UhuAsCSRsWFgJPOVhTVsmBK4D7vAL
LQAuUUAr3JlPSLEfIyTGuOvii7++Eh6/Pg==
`protect end_protected
