-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
jJa8nkYVYEgDXKKafq753LC+pFWhZhLXQdnHn9Y8brwYUqnTFotdVT0P6gdfOFjb4JFnjnz6smzq
S0MP0SO70SAhwAVG5vHwLl93PIGVtl+M+lheEVIlM6SAxMfMuNB3hqMoZPvdQUcF7B3aNTSgIhhV
bJ96x3ihHb5cFqmMtZqEdZL2fIE20dHWAS9n8PMSK4VkCh0X5toVKqygeKn9opFkn8FaMJ8tpaEY
J2cX8mcNsjCbYTMQtUm6tdr5D5Dpq3WxqonHy5vTKG/rU07XqOlv6xPqfHT8YPsyWhgd+degCflt
uP9gsVlvJIqKjD54XS4nR13KEqEMA0zPD6Q1XQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6224)
`protect data_block
WMwpvdgoKDQrmLT5CP2JC8Ms0auHnA/8VnCpi2RZ7keI0hXWfSb35Wqs7dS+ddhPl/rk3/xYVKOw
eC9op4KijPlLaoFjhPOqQ4+9t93Uq2y+ov4+H7NUwIahn/9iUK+YqOPtu+/r4/UgYNqmUlKlJ+kR
boqybmRogrkVd3Si+dSojLz4hXs13aT2C8g+pnlHk+cHyLG6uhbGztv+jymSuiphqVJFdMUuivLX
JR6BBTFtYbdKq21kRwDXv/XWUBx5sokzoRvdD4hnzm94+tH+dddRG4vuRvsGzyDsIEB2oYJQGKu/
/S66tXWGhHlwrhc2Is9mUvnFr29vwpXXmO8ZvQm9RZndlll2lfUkTzXGEG3W0v+4LLqW/hyeTl7Q
7vcDUDTLCMEe53LUgNBaLN/PNK1BfSpz6z3OrKhy/44AX8/HUXHQ0zzu/DO8RVGmNtMINoWMK/vx
7mbHshD5acVTQ6egag2h8Nz7uS1qpEhDNMdmlT1Uy2gtNvxEXGGY1tbk606bwa2N/uDc2YeVDH2m
a9/0umAQODbr2IEZLiCg/G3IjMYMfAkef8qn/M5hr8JJ96R5b9IYnKPWvdY5OT2q1PMiZAoiruy2
vhfpj+jI3jaSg1x+nwbPFS/8Bu3IoWNW1AeuK46WinLPMWLL9DuB8ydUCgVbw9NGlj/HBfB3ECIw
b0rNRpvKaxkQF1F/iD7y7vD3RLDlA9xC3HIhTP2jZXeMRS0i/bbl7JOQ0wsU+acmUT4YetmyqKu7
NNMmOPsHWsp6PBzizT6ukMDCWKKajGsgpEuG6EWzuGLHWvukXW6oz2+hRO0AL/55Bt6ulqnM2elk
pF1dCw26XXvfhWtz86vgMYKU3uXxq3Lsx5K1Bf+k+Rw+Ezz8wwtCUFaeBPKKSS2n9VXsKqOCE+ra
OMc4K4AAvMFEFrUevule5swAzP7WYR7aTh2wRj7hd4Brt/jnkkxmUVm8TQTX8NK3bXpu3xM8PfQi
sgjHd0wt3jbugGw1Bvf1B2RT65kNkMk+yunb0Q6PjmkLjOSzR4hzhK0ImGi8ZCOJlK65zXBPoQfh
oJoSYNiumr3/56SDIH5LhN2YMFstZwHzPBGXcrc69JPu5Mk1oPHP4M//OkJjAMcN6m/SxsayYn5X
BgKUmkcPkRmZqiKzs2ioQLhRhXfYIFdBui8QS6yo2ft8vEmvBWlf6EveA1rfCLuqtn9OxyzyJjXb
vM5h85kCHiN9ddXVyLiHdIKWEx/rloP03OdQFsgatQ9s/fbVatAiPzmoEEMAqe5jsuE3NLeES7zr
mR4dQuehah2G2SnPzvH9813vD4ErHF+zF76dvB6nkyyEJ9FLq+S8QfhbzldeWNHol00HxpBon5vi
xSi+CHj1Mx05QXbRDWFc9uHZ6BcHOYVZ+IO0IB69b4Et44IvLLyvN/6I1QjQ14mzL1wPnx3+cc5B
QEwqQ/4INHPhK7cQdPjjgsPU+8TnjQZ0HijoY0O9Z8ORBzFblvbXv6+XcxdvCs7i0BpxoeRdaaCf
9h6pGsKSGRH45Af0BwBRSZK5P2Pn6Ld6te49P+p/X2lmsDqPrj/WsK0wVlcXroyzb0xrS+a7eKwd
lGoctJvLosba01KrkvKYQpYXe6yLMhVifD5Zyc0E1w3F/fp5CBl/e3wa3p0YOQUAy+q1Co0imeb8
ap1MNXkeoYzq4MA/SqTtOJVvWy97WsPqDMBkhIicb2ot+Wkw66qUsv7IHijlM1AmiUZPLvV8+EpO
FRjFlt5HjImQ1qfx6E4TkbXY82pe/V+i79840+//KvM+bBths77xyl10IxhMHMS0l7t4Kt+Hp9cx
riVV3xh2sJYacwSOboGmQ6e3OvkcOePwlUKFe2oMKGM7TxERGxx5vii+TBxmhQCZwDKe3kLuKo2K
5I9Y+kudoQL6K/dyTb2UCppeSGBJ4J/nEYNYZwpD4NNh5jjzezdgNLCL5eWWiPiiwRH4px5IsN9e
GbUfuIhKZAYdLAHNBV5DW7o214QA8C9mmDzMf2G7gNHeslRL1cDBQX919F6xZjtm1M1dj4+NSgDf
bf3ikWV3HlZXa33eRwiqFEGOuoyossvnfEmwEi1VcAzLuadTDqJIXy92A7DU1j4KNJf0ySpzOyl6
4lT42oYCIJWu7KQ+IKvTDdwTZnU1UECNvjImnCIOjCX6kusS9YBw9VmwM4bozOZpYaYgq1C9hS9q
rar2s9srosNkFdwXI9rgKuaH2lF5htB5vJjPcFnI12xdSSvc3ZQuj6zg3zV+OB0yC1/GtnOSa3yr
mubeWj+iVtGqsl4IRngxnK95R2owuUsOsyajNhnCCRYBTi61n7NtZRm/CS0XkhgDohpZApXTY0+B
2xf78TemVdFDc6UHfM0z+tLzvpf4isuNI9rAb99zIqxyf67E+DFC6TE6Gr5yP6NdIMsDfLl5cxIC
1d1d7MeqixCVjnCh5DJR/uiVH7jOIYCNX/5QCxqhKusyugUYUS61bs56w0PgkcFrexu3a5fB1c/A
GlgrwcRBZGK9G+mHD35GCqm0RGVp0xJAdoMCqp7rBnfvDnS9YrK46EVU20ejtRdSrsrHDTEitmln
11dcEr8CKHoG5rfOnBsPyY2PVryrPBBaUemWfdVV+vZxq3G3ehWE0qJRZ6BF781ApGwDbKaWj55c
RLnCxJyJ+DmqC7/NuGL/ikY0ZBflXl+jdT6gHZiysFambksRF/rfJyMOiD0DQSuxiuVfuoETB17a
pLRZDP+LZ5Cb/RVq1YPyg325k/WcS/vdCRbFC9XCccXOsrFq/ghNVHrVYgmxJuJPF26AFCxPtwQi
2c4IR9X+qBs1542otTs/iqIKia7ya0GD/NZjZyXpn98gqffpzr65tTDRGN/NqJ8NK8c0RqPpBlJm
GCHdZgKxi3RemVerS7suLlZ2ias0nBLY0pJSDK0e6Dc3kp+uaBM1+ljQ0SFjdr5vQruud+i2s13e
CphtsQqONGA5I68YLKOWpRQd5pNicm7bvZUYoTuw/m8HbkZQhBRMr+/dMjHhWn9tep9ZkJRnB/fu
mb/I87spBNaiF/JLLF+aNsm5o9MdU4My95kGJcxdb8n1i5+/7Ow52PX5BsgDgHtWbkqyU0qW+o2Q
J1rFTdK3qLOOpRmX4aLFKL5J6yWlZrkunDBnBnlb+gwqeX2tpYLs0ui5fLgfYcbmf3gFcg0FbEsz
MU+Z94bPwszZxUhQ7JLREFpBPzZJWvimnwgtN/3rr8O7LKfu6ZWHgAEsDMcDtXEPSoeaheKa+ab4
kqyfZJau9Rr79rCzhzBxZhcxR37lzKSVEnpN61wRHcSUMRpimT9JXEdZsHEdn3GckhSwN3vPdkYg
GGoeZf8S6dC38gIN68HwxZavfw8l9za+XLaDpTke6A5eu+DIo6Tj1ys3Ir0IV28hzMMydiWHy6IZ
RIVyS2fBxOW40ikxZHi2VC3XnBQ9qJe7wzWnPSiNyL/NokVzdC7Nqb5SW+tscQ6bpShlWVaoY6C0
K9S0lZ9DmXQNn7Y0rve/ZGSb5doXFCuc9TBnT4xeScVnI+u3Le7iwQ9eF4qLIdSpb/l34OLd2vup
8LubsEVp2PoIMbvgzvAUMAFcdAJFzpZympaLRbiJaOjZf7eDPK/9Xrbl/krXtqLqYWD3BsjtoOYv
FXvd0UG/S79KWzEz8C2s7Z+5Ed8wc9lkfRNMuyULhE7t9aAe6aJj84rfkN8vHvny1xsQur+ZD1cx
fjN89oIY+mdBY4HkiitckvG/JmqFa7UA9Z8ht+enMpiaBfbMNaZMajDSM+fFG3VQbxGjSJAwjzD1
uEHWeI2N119SdW3VzhRKZu9KBV+H7otakR+RThmwy0ceGxdaFNs94fATyTw9pd69iZyEnsf2gG5x
kkl1LrZV7SHYCGgY2wi5yvxtbMKK74y6wu6kEKOgrhEKdkxm/4B+CPAIEMrpmd1rRRp4kkVRGTrN
JU/u+fCMytAdAs5x+L+56ckTXxYbxRlqYLol6C0Yd5HRkM+KKk4aIThK7GvTf1CLH5masi2tisYm
kkZus1Rijd4+g66/LRZGW8IS+VOEjD8EjAuYBka7QaMQ70QyLMeFSmdcV3SSDpraxt+kz/D/0aBh
hUiAQdk3LCkhOe/54gyWHQjcJbKePKbSlXm/YhVf1bLT65UMQskowOrdswEQnFzxML79ypA8rSgA
iIZFGHN6X1zBwUbU84R8Y4KJSfNxnUdvQHdPl9inFP1kMy8MiJzoJLaTnKyXHuK0P8ixVXqI6cSR
7pFZW01qmy7f0pyM/9Wn9qs7uXnOnubPi1aU0tkfstajbK4eSxa6I+wFkZIpfhVyvC+fgCHOVOAv
9Rj3ek8vUfu6PIFA5ilMpECBqVJ1OJGRupWrpyLMnvDhtbxv3LQdPLwD3gW1SHvBsMjWPG1KGvuf
slbvQkINPY/MO7WRD/D3kx8GxhSdry+IUsOG0djAGafL3dRF9pDGL5gSMoLAXfW42T8z5AFUa2jI
Z592DDFxkwieRaH+HbOFARtWPuRo4jvmxE2FsRU/p2ddFh/0/gFBx9Ec/snJSmoVRbod3spEt39Q
hGpuAVk7wxEvMRvKHAVaYLCfTzZfJH+NjOH5/p5Q6K991UbqxUmTGltT8panaRH0H2b9T+HJk0Jc
y6CnVafdRcGu9VSCj/IexSn/3BZWa23/pQdyUb5F0gNx3iNLyvtLdAlUjT3nCT6eH9P46Tvr65Tk
vB6zzS8/mHoCN+dH9wRE1cwqLgdVx9YP+QqW+Fs9KysciTOOUhL6pK4tdcQxUl/N9EqaoM6kqizG
RyufKahQrj2IesYTm5vN+DBYp/gQc0zk+uGEpN4V8r2/QtuYBS9+rFPNIUPHYvvbaoBB0O33C3si
h49vQNTUWrZbgaLalFJwLVCdS5BLiQ2yFDVkMdl36cL2mdnuZPVRWFJukPPYH3yZzLZGwSBe5lV9
+4FvkGt2IDxovt6LC4hXfKYozeLURyqnMeb1ULmjTMMQHy7xOfAYGpydevbYGMEltGTfz8/0KJ9d
zebgQIOnUXS/oeg0gzrpqumbY8U81ae+wv5MmezuvAkhtfzGJdmGDi8x5VMNOhLt6hpi3QK7O2jC
+1axrygYK3ouYDJT96KtLH4+qmX65yuLfzN1fppqukR/1gT3UchN3j672WM6HDHzLMdRI6/hM9NK
qpP5QDPakVwT2sPWtU1elcLrGxOZlYZGDLnqRLF93EJbsBUliLk9CZauJSeGBJLmJQMhdDa0c7nK
A+7SnnzDXMg3mWXUPA28CbvshJXddJyiEqTTHXQyWXwlPtCwRxYUI6VyZ1KWBlTzwnZeF2mGXywJ
DskhS7/5DTiallM5Opf+XpeZPabcUoVM/t8ihMdJnevcbhztIQqnkKi0Ta7vXFuYgT24cNRoFVJr
RVPg/0GJneDLtllhQKlGmPoEUeJr04OWEVuKNYEvhBmXXsRFn7Zjo+cckD3Ien4ekWg4EB2lEOgE
h8B03m7TFfkzdKItckLM4Ira8QIHoZvQiMHNV9wuhU+0+hm3zF0uIS+UWLOmAEnGP5I1Wxpyvp8n
RoU2xzHfptWkLsmp9xXBebcJ2GKHrJPrKLAtRlv/OSecMsfJpmNMZox4btD1ljgC8iaSg4UQMHGx
Ac9BEU8i7GTnPy0TP40ku3Ne/GUOH4zp/XZwthpelywUUVYoW8N9JtokycmHj5m4PJMVBKJxD7Rt
6wr7ocExErJZh6mC1m5qywFrHiDLyWi91vbhwhuf0ia586waDCFqGEax69A4AnpR4joUg6r8KOMy
NyWmlSfIV2SRA5FNPkieXMYzGNkcY49xTnS9DhrcLEhD4/N6PQI6LTYau2HOwySnTN5atcE/1hph
O6Cn+ImAUM0slOVu9nOSewErRWvB5pPt4nlOHxuHJS2EBaCbIVUkdpDY6NUatesPPL9gsMsA8X5b
mlSPg7KZaZaw0hRjd/c+IPwqaAsbHZaOnDQNCSY9we3TDeALcPnJ0klADIFbCXUxppgRufuivjWS
pWTP2XSE7pGuhyx2e/HBqWDn501M03g3hhEAjHBgaStT9r1pqUuQehnlVUsMfRQ94MGqTZ2/Reu6
oW36PpRVE59KoeelrrYAAErP80zT84csVTesTMuhkQSc9t2TZQjxaGUa5ILMBhqyLZUkrQjkwUvs
7/wR4HTKiqkciFhhyKLtFOsQ8bNBWNfS7pDQRapKd8fBYBQeIwR+Qk5ZDxNlIrMYBvBxyrASRDRm
5jVYPuXLfG2LtbeFDzwd1Tg4rk0MQuCEVHHLyur8wPH9ZlM7n3qPBddV7EfY1E6PhcYpA9bFc7E1
zFk7Nldw+onhJLf7wPMKwYyliR99J3qsHS7P3wg7Tr/b2LLuCLFs5unZMsIJX7I+N9Dx0zHIUNFt
JYtWte3o89AofBOYJG6NVkOUPt5kbMpYZfh+20ZeIDVHRiMjckjiSj9NdUmGBB7RNUzp0CPP7Ese
iwLqDTYmi1IkPujvNqlUl43B7rFHDHfj7xjsFvXPVwfJ8UVYZMjhEd7Q8Xv340WFlbCo5DTvTFhw
JokYdSicscQXcKwJvJTyfsPEPcrLu6Ljf1zl6zt5EQ93psqcs3dOQEqRSve6qyqOrd3x33Gklfpn
5iHJdBE2LcfgaIisQJHLio3p7koqcz6g4/wHqYDgebhnwYZIsfmO8RxCp6LsQZ27tsLGZPgJmtcO
HpJredeNcxuLKKyZab2pmkpoSWXq8U/uIQgsxJcpzQROyarTG5v3Xcq0/E5Qo5S9c3EN+wVasScG
WQIcv/I3HpAIT4zYRI55Kf+geD2tGiA6KFwMFVafeWpXWxNE9klYasSZtuzgPO1OReBT8+/zHUjj
lOKfv/THB6R/FGWKnCZhg8x4hvS6ZUhGlYQq+oXNQZjth+I+JWNeuxI5UlhTu6v5i5o8H8Bsu2LL
EvwPVlDewgBFCUYfFuoux2qQpJ30efggrdUzC6rnpnL/svKpjFMuGL7yIADiOJkMdtRjEZJeZFRt
gLs0OgDsZwPbciD3ldnn6x+0An+5UqcCV1V5kzYrzN81Js9cAW4Mt2u5MZjlZguO0N6EuOCfZmeR
F68Zs5IJFnvBGadWQZxDAHf2mEBmeOCxd/VghdwCdmixV3q8KxN1EXVTlawfmHqDF0WEw6s0P34d
caow0F5YIuF2WRF0Jt26arBbAeuSyGN4JZV3PGtY3/NzcbfzktrgQx8raSQvCPmMCq0f3TZt2EPI
ZvZahCv4E4psiO/pZKAH4t2jwf3QduDy6wmyOxJ2Mc1RKYQQXjzwEtiZfvZYiBMzgCew/qxQ1D5A
AZgDZjqMGd2pUlftMYEoKGV7nef8e9bnya4EMJqPfg0GxcBPi8dF5KK/sdoew3sKmwDvZEPXdzZV
Be3ulkfVOE35184K9880e5FkoMYLI6/x4sX7DeEfBmSdflSEMIaP7KoTjycLGvf7ayWK3jTTAuyW
E0j/wUARBJgQNvNWv3p7dAzNH/J9VorghN0zt2nAWfOejyyqJMWOUiNgsP5oKqQmw5F/ss/URj74
a74NstCeBwloQKfzoy7FHv1xRaWsiHXe5qLwOKXv+ESacU82/mLeUFRmQA+08cKghpJu8WIlXlSO
+VXDXn2GngBdtuRZ3SVVpJFfQdR5RshYMJb9XdYH9BZtvZ24VCIEsL3/gLGyL3/GxmSvL39rauLW
Lnwc8zFc7Nmc+Bz27/6IAa3tPoAxi474Js1vax/t5ZMtdqyvbaa1PAZIrYZpgSI0ODlAJy+fg3XQ
rBIWJTiEMqhAPPtRME7TgCR24yEvRdtn9naPP72ZH440hxyXhSopVwUEbwOCoXSk8YlCxNScr+f+
n4MpAVn1uQAsM/x5F1xPCmkx50ABna260ZRYlGbCYlnv4Qt3htasqK36ITtxL7V8fc6gInEpUZDe
GFpjIgv3gNK++MAqppi3ACxC8oPFt7N2XNEcYS84LiuGYeh4sb7LGlSTKyVGMvfthO01gwTNEr+o
/gPJLZSDuf8r/wQNsBGPSEZMgrAeJWB7iV8G/tBh/Ky6nYGuf0hvDsAWMNreL2Yb9nj22MGqJY16
vaN9VJUDYsbeRINlKVyhgsP79hFcmIpH3LQ/vCC0fvUBQ9vKVstZPSC6SFIq8TrgP4FpOTwgu7dT
FAMQtQTo2Thp5cHLDCNunchFbwTlIz/v8PWwaIIzBlLJeJmSe/tbLqIkRqdsFLlMxKpCOjjZYc+r
VcW8nlKrVzCwI/9m0ZzINpVMneQ3udHg0/NUJ7t6pZTUYLkC0lL8GnuKdUbkrsiEgZhYCxwshc3X
I79N7Lyop90Zpeo=
`protect end_protected
