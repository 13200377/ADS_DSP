-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
KiYRgi2RcRFYrFup31QWlZ1d12q/ZhisbbXr+UbIW2C7lyegQQyIAZo8+FZe19ZTDOkIBiR7AfeF
LYHT+dqBsIBjxoBcYPF82lfZ5F8YpGy287y8xHSW61UOXaJF0kD/6yd9fIgyzmn7GuTtDzswODjg
7/bx78oSEPaHiCr8bynfywlU4uzXsKFtq+SzRHmZl7s0fnTuMkuIwm7Mc+ePfNlWQmdw/r+OCjwl
fbbzePxW5T3mFo7adZ3tnvmrOo+qjkskq/prP30SPC46lx/0I4Kcd8R12y3zw3cS1rrO/uNyEoqF
zt1pqC2GX5F1xH49OwMAvzT4r5w8gKrbepw6kA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1728)
`protect data_block
tUtjX4rnoQlEvYHgbcqjb+1f0Ys5aY9aKfTPGZI0pOEVgkwPwojfzBaILa2RjAKzf0w0UHyM7z61
hT4Ev9pShYbQnhwzdMKE7e5zy9E33ojgx/Bu6lO3MYacN+R3FP1AJG4S1vF0uSkSZ6Ac13xNUkh4
M/G0wI52KH/XbFAM5OZ34FGVPGsu8ir/RKlwE20xaKJXZv4j2fADXuUV0WGjGNqedjJyrmUpqCxX
8aLxDmkpl5ldVEtGAd5k21V69r2DvRChU8LWI28fHeqz4z/kZWrBiUkADfqDgIVx4yKq/HEP66kr
VPXF8sJXKSLN0eOEv+5JqLm2oLY1vSy8mT8ovPIBUp2b4ioJvM+RJUfkfld09mM2Dq5y9/ZvxGOT
WduzmDrJQsLw0aPOHPAFjOtfCOmb1CM7Y6uOKwCk2r7RdBgAi7riQDxPR9MKySEYqDiirtxu0OAA
63qAHZPqN0IAQ4yK2fTWWjW3xkrYEutS5ZX6NbCuGM7nmW4mxrxJfmaLdPWrHQPvkTbOu9z1EAYd
XID0xygJXdw+vSMjH98mQBfhOL1cfftjyDxAaWRbIEeJTGQc8C5V8M6cbvxqaecSV5XgcshC1pyn
MyGo6UuviLpKh7tHdtPnLeZ/gz5rz9qq0qeYseto3bxMBZ0OmuHqpXjwJqig+QpGIW+SQCrGVwf9
PVxASdx0n8pJqktCnILuGavS20W7w2mafpIb1uqzK/q7Mz+DoWo9HiPB5o4eQVz1G7nGILg2uPsG
mI49RI2QccPzRGhfhpMQkhJyQH9nvRVzKRMCIVbmTUi+L01CxuAwosobTIrPbeM5qWSfb9d2dF4Q
AOZKTGUVZjjZZgAeYoK7eETHU5Nv16W1aHVwDPhpY10coHrMx4rPxo1xw8yQvkO8FS8PaO5yGCCS
VCqeX8SlKMQr0p4cDfk7TupIDV9tQA0fko5hy19cWt58AEG4lbI7FweWS7L9dlSeYNh4Nfchwa9t
vior9nbcqAJIEccRYDxcMINOPAB5232FmtCyJR81uUdb6Iv8PHLPc0vgibGfqgsKwl27PiFe7k4L
gR7mrWSeWA1ZKZWcSODuLi4qm74X9D7xO6AM1Ci2I2RPU10KbE0M5rY2hTABmISN/V2k6xOmGcfT
fgeJEgjF2hxp3O6hf/tMcS7F+YScihaqV3Zq1YqFwQ6KO8Md8UmzVb8KTqxNqi88NeM6a5wYLCAS
U8tTcMzuzPb02hEGfEMIUanxkHFNOwTxj0rw6zyJPbjLxOVFhSyDXmMlsNXqZN1WjWO5v0R1pg65
3CIt2hfLwPJW6uPMRm2MbF+uS5tEtV0HqbwH2qDC6tn/WCt7d2WwuZ+SGGNSiBLbMlbkd3YSTZiV
n3TTjEiTap4NCOpEMaqmxk+UWIR87pJIVd4tJLlRW27qj0ZAgUM2KDrOaz8NPIGC7wjQmFHTgctE
GoRChpYXylkKMh8F/Rt+gTh58dDFQLGYJpmoWZ/6lF9h2LC8SJMaIfxKEMirc2yGfwRqAYJH0Dyg
54hIV9STR3vu2g4zkLHwGY7Qxr04IilGLou5HHeH9ik/nch0SWiJgB1NBlJ2DismhPcfiMSKyavM
ly9oKfRITzvnJMhzUZVt3ACMrlOa+0IgZ3VZEz3njZchIEIN+Dq9/Wdxsn2nnlMnCvHJFmSwXd7a
uhzFmnawU4yZZaFVOko8cLmwBWPbm5AZl3Ty6Kt1SQZLJ74jICn4ZQM4eL1FoxuCWsY+LDmP3bTC
bJQBPPd0agd2WaltfyQeL6TC9T4TwPY+zjlvDr9JfzQ2UnFCnGtyUEhPUdofmTFEczGlicmsHvRV
NDUi8Nnaq1H6CKYF/Ibb8rStG2er6RN43/QUUVD9JW3ZGpT3iprDE3SH9NURgbTkg8Z+AwvPWwM5
BkYs6VtzUk9jp5BZ/DyPfy76r2+gU0D4B5/ULsJm9eS9A4e0KT8MBNSByFd4EiWKMoVGgQfu1SuG
YUnO8VUUeftM+n0Ys0QWpDn8YZnI9BABD8OTnopV7E8nTxs/wa4vF191qs3SkxN3VrpMMUlDe9R6
z142Cl8aP411mUsVfZrZ1K0wqqi1hq3w2DLLOpsaOxdb6y3xC/udlUXlFmbm/WIWT7PLU1jtiKLW
8yyWhqVS5daY1OocXwlx7X7aY4RLLpEZt9/kdKllwcAfw6EVveJ16jut3hrk4tjqTQQLhSJlojc2
yiowDBqt21fL1V8+8d3qvjfjLPezApKdakMVtg5AQK0dDzhVJZXYGxHkA5MyFhV9txIWOAm962gB
noAJNEa8mGJZGCYO3E4MXesr
`protect end_protected
