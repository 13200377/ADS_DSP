-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
w8VzR8QSu9FsK+Mju3846e5eo3kSTseZ4hAYcqDBmlQDFNldNnQSIDYiD0W88A5YmNGmViO4qbfA
GZr7jThDbKaXp7q9LcbOjD9iRW5bf6FqCGSHK1S6PW1Wl3caC8k0p2cYsdGQnoG7vHRfz9GQqn5K
yWvLdNpT+pYahPGbI39PSjVm90kUltOnpvPHY94doEI/wrDVUya9L1EeBviyO+Xxrog80KixHCtG
5wCMWDEQE9h9ydSQXqooya6AGh5KZzBYPOV+ROAu+w3XyEaczxbv55ngqpc3U7EuG+Z7YSdJOBTb
3R0rkEaqLUhfo5ABmjMqR9Y1rKwWXkG/Vij7CA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4816)
`protect data_block
ZbeL5EyQWmk35Zsl+5pQkwT8MSF2ibKG/TRtqUTUhw2h3SfnwVXZeqHzrSpiOLR1gzTIG9ZjbBIr
ahr0uz2hVQiuihs+IYLz268dAFkdAKQx5bkzlsmulR/w+wvfAnDq7T20jqpelfWB86G3DUWOhk9n
Sr3H7krsNysPBxzEmYIXhUWgodkT6CsJRR36+mu0bUxJd8HaXxM5wOXnMmQ4SG2fzLbQ5wgB+srM
0HlmBRxaXNn3yeD9POJJjtTAhNTxQOygo6sBlpGAFd+ZpwwVR9kNP+fptz6t0qKs44moHa65audK
XTPflkJV6Y57u3sinnMSXAAlKmckCBNT86+HAgqhFJwudgIriJuGabbu9rZxzzWnOyVgt2aD2meT
S4GTB0t7g9JSQO+wPBPEtNDYIZ7qcoUiAL+m7Ia0yiEQPk6lA+fLtnBK/SVem68MmSYVZh4af12A
Nt1m180H4f3GcbbcwCfyh5fjrGQk1RVXzY3BYH7g35/4gbt6CvCciwiJbXNVXgiqftA6vvmjzmWG
CCgT31TkJfuA8aRAqDYcaaavVPc8d5P5v3pSSkiEdSmDaE5wSYpV7d8aBB3fM4dDvJrl2a89bRse
wdZ+rTg2Yky4uc3kHpJoTXEs9dsIAqGuZhVHGWMaQYpReZLhaxDtoNCkgVsKZAs/zIrvMuhcT1Ga
RuGkqzpzHSqgXNLFy+NuicByO1aHoYA3lBB8G/ixeOElVv+rZhqm+tzFXU7CY3fJbdn8L4VB953z
BMfK3C79u/m7xDhJIrmY/EC+rbZJP8i40fG0dhyZdhbc8nKZEYs7OpVYvtnoLyoxcKB9J0g6X9iW
Rhyx9lgSuCogdYblhuJNGBsHddCeRvTX4y2tTjEKp5tqye7CWhlaRDSRtspTURVBHOt6ygslUBRt
wkfg75KcR/RTZ5CCb1NUgQ54NoBEBiPhsB3g5Hj9Wvf6NC2GE9s/lWL5IDz+0t/CuT5KCR9i2Ato
rtKxTzxDFMpOOnN4t2JOZ+DPUTuvq4N0oCVq8BfQ6m5ogli1+zWHyzuebtoFzZ514kLI03zj0ehd
vUIcH3qyAaykM6LCITdcs/INN+a8uQR7MmVdk7yhxGDE6hiYzJj0NcpoMHS1ScOMsD4a559FdW/B
OmOJ7gHCGObw30YsAc407FIPDLl9YG9My9MxYFUZVpVM2v/VzKgaCoAGjHEO+XxyJ7BrvAKWHMWw
fFOWqoAyRYMY3E90+n6hFv7/8MXepgKxvi4nSP34ZmuUOap4XELP5GhCL5nquQFLBa4lEc8mr3oV
cUA7eRpjClyj+tS6CANBmJjrDvHQTH4TV1t31TtN17LOQSoTLL9xKhcz7DDzerfSfbCU5gfOji+W
u0aD0+1e3PX2BvaAKJF05nX/MmVHgpk1EJHlYxFgsSOvYmTdp+liINGxSuXkAT24HC1OdXVnp1at
abKXKL5fn5M2LQcam33084vTUegntjfTVY7oDE2xk6HuE+fcPyTinzA6dj20meqGwDZsccxMqlBB
w0hm+P00zdbTGf7abnr4LRdrTkyuD0MDo6JKPt4nOTg79NVVKQEcj45OzBDVRH4s1RRY9WNqwfpH
jAFx6X2Yx+IbkMOPPxxGNaMOYXhPgbuCJP2j8cve3YW97u0bQ5i7v467dGPLvgWCpKHef93ziAEL
5zDc475czsJEzKWJ+/lWJuY10GYA5IFGO783pQhv9vE3kY8d79RP6cjQ0XA6vNfk8Iv/bsHiwndc
1yoJZrMS794qKIf3KJMgQA0dTKaCQVuXQwlePFkaL9A8OLIte8vcGZWeYRZ1D1CR3X46qc9bamob
z+4XfSvBRGK7ESlJltib1SR44Lk3WS4oPnn+8DI0Be7AwTkm+/oRBjVwbGMIE082dk6Y1pBxxcUi
v5MgbgikXOhHzEGxOKc3XEQxZ9B1thr8k1RbWVhSoF6QAG0sCxuaI+t17BpbLyMaQH1ZTZSVzLVb
W3/Oe8G3E9DmVFckl6Qojhq9ExkQGkNeT25Rkqgd4MJMf+4Tei41hnwISIfDSJTtqHGWHzoMJn6T
MZfz/zJKOuhh00C9PJz4JfPIhOvupvjI7sxPRIyM+cjdyPt3nzpldklDzhP3DL/hP2kTSisGrR5Y
vf8zZ+wJXZ3vZZByAMSwzo0ZqryqkEsqpwQF5i4D1d8crYISb/Zlf+dWraBPtHLWY8jleNSkTaxW
jlyU+jiyU0brnbAslt1+qj9GL42NBrPfU8xQu03zlGoQSUnYmQ01A5Xli/WqFy4+NlhnA9fzx8WT
9Q3a52BKEcuw+hlQTZCXFvbamZpPr8eTNBso8PW68/ubSpTFwuZpzIBgbc+Wh98nMIeHbXCRT07J
R5iBlhlnBMZICyHmDJ5RhXCCpPkPVz2sfwH/Aj6eqPuZYM8wjXTdZFAKjtJPbeC3stlaxnF7t3li
W2+CK4oVxu8+97eK2Wd56slrBI1j0D4Iw7HyzIcyiNzr/4sOnckrYEG9DB+vsUHOQ7UU0jlTbEPc
B/4js8hLwSkW+8Fcq1sI/Uhlm35ca6RT3sqGequMzsaCfbBGtK31/KldelArXeQve1pWdVJdGzrn
moRjdIFoMHz0BA3Zw5oGcQQ3tiA6WkCXQwEK5ZxHjCks/siLG+E99bT6DrsLRtOHa7QNEvtkW7AD
5hp/oOIzrAhSGlwFBiKqUoisvjcJUOGgQUutCrh1gBsmmT8nWAiXAKMIFVtdSUQJ6RLoVbf0nlbP
+X8gfEOZDEHvWmBLmSWyz78XwUbn8QyJuedFhFTWP8srvsGsTwnq3Dige6XzwmbCplIoYI37XXsW
jBalMJ85CDYURjeOqewLWPk6dg/M2mqFYMswPZE9pWapEvh3MQPGZaHSY0k+DXGP6BMyEsXq8vfp
hBo4tr92ZsXIg1Xc9ylSYMZnwctmPle114h83IvaxvL0BwHMd1CvUaMyAyu4ntrLYFFNeXIKRILg
qx2GCvlpYM4gkrfpPB3JhBR979qy5Hl6iYkcn4hhSbUolA24XNTnzYCbj4KowSmCKYeo8VYm+m/4
TXVyx/dUBjK15IF+DowxcTe9RMnn182ZzVHJjYv39uuNoWdwW+VgTVN5Zp450JSV5ZcMFJNSnA+b
u+tyDAekUTOD7d5ME+aJYzPIb0JRIN7IpAKLCXAO7wIMl+o2HMaxOwMftZ3CPNbcojW/3j4MFUcT
zCUFZc/VtEfjI6SVcK0TzCzag9stAPP4xzJcRefTgCTJ2+Cyw1du3dQq+/owmTf3E/ce1sz1EqSD
qxjF93q+F6GykQ9D5gZ5qhtLeoH88V4EErDhyTgTUOWwQCzsE+2B3jRl8rC4q3+mUqZQ0kvUe7IK
5lVeYbCgTj3qxGYnjYDQIY+sqi8qWiZIH87bySLO/kyJ75K3pNHa3yxfejJldqBIK4SRULX+EhlE
G3lAneJ/akQAIkxavWm3YposA20DRNuQkEfznAFrzyiiEbrA1hDcj28XufJyzq+P3vZyc6H2Yrlg
AkXSc3ZSFNy6DNY+e3EjUriIzeRBDcn+zbH/21odB5hTEQBhUjLdFd7t6o7gECSPLV8dCgEpjmQC
QZtCZdJwFnXhElWZQHHnsnJqDkZb2mWRTfVTAUWw8+x1PlJ41IhxrubE8lc/VMChDCWvmx/5QHyn
+IQu+XRwl2AlT64rmyly1yiR7BsvE1IN8MpzmnW+wt11y3FDuveqOemjq0+ffps4X4sKQjrJ3LnV
VNGjELJuABWWH67JDp4i759NuI8HZyGUHspK9slTCFl1fLxuRdVB2BsU0SrPzhabcykwh8AVqTkV
AN2wNZETHDuXqWenmnJLbj2fsaUFY4A4zxahchRTqdL9Wfgq7ZGtilGFUbnsDcefNP3lt8MtqzLp
WObyzhV9WpWrILEhYlOlf9GBxrj7sEmfjJfu1MAL+V5LhjgtW0p18iZxKWRIEtQGWSLP/SBc/08t
VNpzPs8Sahq98niAoSkWGlamoqi16bY7GRIxDTlipcgZkTXwqyDEunvKXx4XA5b9eSmSixZ1VAQ1
1aJKrIVOyonLwYM8Jj+mIirJDNaddXSBKhKvmQVc6kMAPROQV/E0cvRdQNSvk9cWoMe7g5O7AtYR
9f/s/GM36aTomll9nQMQdQ1xF2F/VdF/nZGn60GGieEGK/HnunV0q6FkYrI/mWZBsex+hDxutUkd
6kY82PJgxbpGmHzNwIOt3Eyt0F6j9SNoEbWmBBZCw9Zah5sXE9zT+RaFepIckgyRuXoD/FMO6aRD
msU5F7ZwVEstQKSKCXrdp4fkufGaUxcEGaZCyV0NUzeInHuWFjteT1f2cu8m6suuVOmac/Xkqcne
zIPMtb+99nqriEKhkTYBR1nVvdQA1UoR4d+CYrTOgVWuhwtKSBm1sAqWc/8/+N3DLggij+hnLdFn
rmkdMsMj90v3TwiklelicPyoNBEnJNeqj/VBChI58AQVphPfP07E917DP9PxSZcqm5xqVQ9wT04e
SGuaxMbwfzsNO4CJRwZB+VSSpiFu9e02ELxPQ7rUt1po0Y0LwWyXHumOSA3b+tnU68KKXQtMBYVU
xyH7fXRKRKrLyaozQLQ3WM/R3qIZK1o6o5IgMxUPyQsFfV3v4JuTBHLdAhaoaT+AcfeJjDh1MzDB
P2OLlNt3zxliIFE1xkzc5yLEEb2+pcsrah/pIoiaj0piIQiggHTHx7bboW1AEGY2q4NEPy1BNYd6
XHO/M9lAJXfmUipqtSMicPcXZt4QMv/vN4LX/IdPsGOcEwj/exuu1aXln3MDLJGTJf+/B91ZDINR
X8ZStGYSeSjdun28NXhxEm3i7JLlsEROI130vv83cscUFdhDasxhrpbvQi0yZlgskiHCw+U+C4mL
JbhOGT24UWaQXB9tMOcxmZwQoLpsFg/l6zJGI+cJIuSAKsCl9rnrNdjjFtpxhKBlIkvlI8+MzRjC
fo6mJaInMLig17a3TvoeUVdTImvxrcLiN7PXjylOTYZAxblGCPkBKna1ehbc9rIKboV808J2NJhs
q3ssftqOiqmMJOzYwIt1rbLHKCNa7qgvp7Q4SbKg2cSc1u1Fl3K6ZJLB3Xymz+pDnrlJ2FCBLedV
Eu9acOca6zyG743CMWbg+cqWb8EkOvipLcf1mPmtSS8a/pmFJAUPjNuLUA05xdwaz0iBXsYBcuPD
CrnO9LD5N8Hm2QRtXwYoPSlFwKjozviOHZbtzg+C2ScR8lwVHJuFweZnmsZld4N2zgAEVHgrNm8K
OSGQsP/cWoYMcz9K6g8hsRJWtF7vdg0DIO5PffsTNlC569SilquK9M3jwYKRfFN2QISKzwNAQ3TG
Ma+rRsVFPumgSV8RruZydQLjHTKaAdYuf46ykkuIktv7ynUSYup2HEfhBB1qrNS88DX4XI0ZSCwo
U3o31+iq+PCT2KPSAiUwvuTnq5bhVLvbvJqNRtmhzq3FQO+MVJ59+TXFkW55UdgkVGoRu8qybnkY
6tBS7VJQDA4SJwx6CjCxtxuWGkxZDv9YaH2ksMKWp/wlrU02wQlKUv3sGyvfnbIT1FLGbxZI7Igk
fhOf4B8sugFYdi9J6GcADcr8tNo/MxBzauw/ymYXWudI2h9NIZaOS/SlmLJzKZWvrsIcFnatLYW+
eANmH4tEgzTIqOO9Ft/y/icIq6td0fls7Wa7tX3TpHNVd4AiZEgsDhWV414qtA/rn26UZburACH8
1Lp16ln/XK4OMsCiYSJKIBGemsN00rYTEJyq8LWTrNGD5Cz4WOyWrWMu4z2bFg3RD0vx9XkJ6ZtU
GX7rN5Tt4sUKVC+kMFYlcL4p3gBHavimkBUzPAYkN4QEZum4ZicDnmQeswOqCHInpVc9+Q3aybSU
yZ/v0Q6CZtdzaiBjRoQt8zO5jhgIAdtT4N+JB3V7RHC2rNqoj+pBuPVeRVPY6rEmEKtY2UA2kJFj
0B5vZzmn8TdSp/CjbgUx81O8BEqTYLLzvILbLauVnAC5uckoMByi+1Ta7cLAYN1ftmTglcndqRG6
1B9/tIQN56iG2hg4w8iVMW+g6zAvHYVefBfPESAr2ohQiKu9/5n55OW/Bd7SNZoYtMJgQu9crYIi
FBfgV7HocNi2n91jei8oExVtXgleWGrVlg1EQAwCM/TfGjE86WwmQ1anjxUpc8ITkCIDFX7qRs4u
ckHkVeUD3tpYFmsvBUHryINCc3ocYI7hLp4U0B75ROFU2ZRsZ8lI60zBMBNd8pA1E2qqORau2b1F
ePyT9opbXjVMgVU/yEmWLmWtPJO+wD70duNcWb8v6/JtjQe37uj02sPJH56RWoTlsd0zdW4+teOT
cs3kkios3yxPwdCcUKnwKEHZrsQ/gugVUb7nysaEx5pHVl/fLe9mZwKja8iU/LBJU++OTJko/MxP
k9H/CLaOwR2Wd+WjHtbJkx2W50c56aYOB/GQ0Q==
`protect end_protected
