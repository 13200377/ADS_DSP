-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rAvFYmcGPkN3KlR28Smf8g4SDVLSX5El4/IWT6/uz2KZLviLHMz6TZJCGEOmPyV4fmsCFI/piT1v
0NfISnjhOHl46mirAg9YfOJl3E+kSggKUyoSd1Ppryhx+mrnbNJzXcHhABtpykMy3jqfZNiChbld
5uIveU/5AtyKq/cFFnbJbtk7L44+LQ0VmMmF2nX8dyrzAPeTN9uT1TTbcHa0ubxRIh+g6UWuALK/
RVh/2iyqQNzD38au1oXSKWSzDK2PEZA+31cjy0cB5i20b/zrmusjprTwKt4KCEWIXKz5eMDK7fim
TON35UOF7lxjxf8O0e4Lzpp+KbPhrOom6ab9rA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13456)
`protect data_block
uMYOFr5GCNPQPMUXtQvJWGsKyiVpidUFK8DjIHq2cBX7hKXcIvH1D7+LJBGuxrvJ33brq+r9LdKJ
UWBmvzd+QcIN38b7yngr69objkxKAiKq23BRZjt8PgidCSzErIiKmvxaW9CVegWGkfLPCU8T51oU
olpdDzZkmPIRkuirDu7FZiwoSYpE3Fq7GwYh0mtqW8PUYADiATwbTAUJzp1R1hCniwlmFrqJ+Dmw
F9phamhKJwf8t4KHeiG2LxrgHSMm+PneacJ23fh2HtUO4QUi41MduEr4QCdzLPgyS+R4jLGXS/rq
RSVjoGrlPjcTKVI1IypBTw7HcdVrau/JHjsuxm3CDdRAnJF838RojEw5/lRghbuBcq/1IpEUJO1h
E1wRmMfofMBs1hbnGKhkyvryKSgNhnh+Hxsn2GRvaNl1Aq9z+i5u2kVE6/pNXskQc9kGetrJTmAx
ywOfxhGGiEW2IZslLOp09gFW3DpllQvvIhJZybZh60RLBJjDNrwyPP5ocrt/SQfyr3zo1UX7kANe
mryiLDT0T0Tq0QyI4BNYjmYP6kChM6mX3QvAU6c+/DGAkcXnGIOg1wEqCNsUxkMuRhgeqckYKv+p
7vUUqEUb8Mf72ZgWPR68oSSS6+boxGmVxod3iDHp5t6i+0bzzjrV36w0CKaWhIpLMU+m4hCp+kw4
kft/vWCr1iIAsQ/URKT9TGNSMU/YL6WhtA+yg4t6hTxj1MF1aOXVPL36+RNarkGd04tPBInhGuYl
RI2K+pG8H6CC4S4HFGYYQju+UWO+NBbWIsufZt9bJURWu9Lge2WTKsB/GgCtZgPeNGc6DHwPdqSr
zxe4b3/IGq4T+o7ZRzXCRRmILtrpizyIRKciSC36aK7GQU3ZP0nXmQ0lerFSW4A7wkygWWPNiKSB
d0NfZ0Ds2pMmxPaz7d2Kj71dMZacKD3M1S2Yj/Gv2nu4IcQKJeM0uMsyNwnENu6vJ9xwIwjCpOHx
5rR9qNC6YPAsILRVujsxo5E3dQAi9Oh5rPQj0qErwE4cfeH08DV2pvKVFBaKgDu3eG4MA7CCVhw3
ANC1sCj3OqypuBfvbHh3deVKve0792KcMY4ZmRZ692aHMDcuF1HyJr8QYKrh2DyVmPObK61W3jyZ
X4qsWRept8+hlheMaPUn/1vfolsXVU3Grr75YZ+Jf+ur3tlz0vcowGERo1Nwu9rsY6X9fKfVK/1B
OpLXz854I7kQjVUZiKqA9ojSYpPhUUO/sx+8ijEMFZGZVf9mzzWi0XkVO4Fh229E76Rfxf8VczGv
LT0IYSk30/qdy6lmpT9qQjRn7sSrRzDvIa060mQ3u9yFPC1ovAe1PVOyzhCFFUjo86+2ZMTEh87I
QGJZIh9xdt1L/4BrRsvJSf4g0KiboqwqOoc7kSJ6zopCMBebW79flASbYTt9XIarBIsQXuQkimyE
dQBBDQOkutfsR4zzQzu2bTrugVnVDYlKNZWFY/buKiPTFSGX5JwHX4z3qp8n3N5N2+wAE3isUrVh
63qT8n8TOTZpa1y+Yso6XFnVexCiBLhxliGOQwQOgiPnlKbaaqRGZwO4aP1FnMP8ah57IuRLjvpl
bgvF7k7Upn71N39jNOBir0RWesFjgYh7pt8Fjku972nhY6XVAZ0rtEhKwP5WFfjl4FRi0HdbcsIR
ysNm/ssJFnVgSRY4gNYUvrda/yw9SW/vOiolg81Eyc7Tw7FU86OjfEIWIT10Um3cHVPSezau/BJu
0+ij+Ot2JL0V8+HpzMoFulpaJZmgMQ5dutmeH8+16L/RM14PhDy/cg3khtL4Tuv82HfMw/beChet
ncSz/9wz0g3alj4mfFiY4KLhZu9emZ+yHuOH1KQFElnS8AZCyv9Klp5xmUDqDAd/Ja8liIBHn4d0
Q2o7aUWMtAQ8HT/OrD9T+Z3dRciQs8C9qLTovzyVhBHhoXeTEM6VS9WhBQcXYcT0U13w0isZrl8R
GJaQfgBHR5XDage8eUG3r6yURza9F0PwHD6AqiNVD5UNiX+Ngbd9vfCTZ/7kL/vPyF+iO7dHXmaz
2t+Tk4JVBEdqdb5CyV7rXFGyAyvKDxVjGiERih5BGm8tOvoTznIvCambtE9W9kA85z/Nek9NOzxL
oZSYL1K09bIORjcSG7EWniIQj6HXSe5e+oQMV6DHFT0JGTV1d1DCgKvb+sbveTYcAvyqZPlCT5KP
544xqYppy7yYOhi+L6dyqG8udYDwVJ/C2r2iYvYTZcgSdiWMcJBbTSoj6aGTEQd2Fr4HmC1Etb9D
klLI0ZGAKqzg7Wzfr18jl52bPA7TXlQ7xwQJoARj3HjnSvo9aRymydOck0Od6iOkNAuNVNAZ2Pjt
PCBLiP+oP8CCygmZ2y2tEtF5HZcqgMeAwQeqo6nMq+sj8MIxt/Jq2mbhrr0zCTa0K3xh0IaU5/Ju
0Qmn/8TiFSuks60OFV5T0GWbxmbJ4Spfbk+WREERutKpZWehXPytZe78qdsh9SLXiK7Pndqz3E6Y
3FMWOf882p/i3dOTn4zlmor09DUiCyWZOcE7lpuTh7M/QTZ1Z6eN4wHDKKLYY+QGQ3oXazmzVtuk
H2qLKtEdQT5ve4LrhKMpnuMKNWaRbkAuhUMwiSISAInme1lqW7hhSjdke3Bj+IF5naFTAvPMAWC8
s2E+1kRK7lxqTskAllw2eTALFLw9mq7auF5jZ8MIG+8YCP/le9SMZiytQodzeWNDMIRidmzFVude
SfGMllGsj89SSxvW0SusiND2NtaS61IiTp26dlZH0aSSmkueGwXoXIzgQN3Nhf+PSR/0jelvDMX3
wsPUNxJlohLL/gKsDfdkOQ2+c/Rv4bmknQlQhL1J/NbYtkhb1ygkem+qmrBAw1CLqsW8/8JlmIZJ
tFi3T4boRpNtoSIsp9py2aFt5cBTwqfQWT9s5KTJ2M3fGDGL9KmjOnlsBzH5Ask2N14jAV/4HLni
bee2heIF3HPTQ7CHhur6bijHPzAyKu4Opj9Crq6xNyZdSIvrhg5BQyF1gsI8aYXj+NznyYVWXxjc
dXBzxOy02FqRcpAs9CA46vs+BI/0RFRHfmRmS4bGMIBbkr4H3WhtHqB1viIYgKBXO0O8M93iJi3J
yGXYlYJ7qtHMkjYYJJ1Y2YDkPBIHGuCUSO7cNvX90vRZARq3+uf6nUb/1TSK8vQuZ6EfQR5KQp6c
+YBF3iDiW8MzdCFHVFXiUg/2Zp++EOtVE5AT4uY3pM43qrwadgUFwjZTMUoFcnvAvGv2FucpHWFx
gLHzilCnnKFVa4+agXBFIdXOScYcdQPw142g9lQWxQRAIJHEZIT5xo6BXcPHMKdnUpA03Rwd72bo
Lzzs7hReS6gP0znCSBLnffD9d33g0Ym9zR5u7LjoigmlXhKzff21MjoBcQRtXSA/7K34pwvbPbj0
hLiBKJDW4h4OGBg6kz7QNta3adeb2h54EMAgVoS4FKxPkI5YN1nlQLs6S5uMg8QFNyxOE0MHA+IC
Adz5+oqunsJMYEVVnfD7l3kOEOLS2xacoZxk8+wjO14MxBIRsc0bNJDI9ZRczhj2K3ZGpRO+8BSg
+Nt+W4PY/1nj4QWr+Frrsxytx+d0DDUCEOURRx6AjTP3hPA3MVhBZd9U6h2msdxJVcWFl5NGikPq
HhXEDr1haDopQjsoF1Loz2iN4pMObTmYacnLxMBIDBXN5rcDEPz3Vl51DBPdlkhzSM1qCObFZPBM
yEnoPno0sZhOAkEt7FOalDaCpmdLtPKprPGe/kB5m1c4J4f25hEu1fNrPY/KzTXtn2jGEF0h8SC8
PfFH+YOt5TBqe9sAGb8+Nu1parZ6JfNMrZVbNgjXNUHzLAr4zlr/oE8tZhCDidF1V2xVxCj/MQVB
0Njx/rngURSCJc0fVQppNt5iv623dHMA65xEyHLxnaHXLeKOVgZMG7q8mFO0Icph2/0engOtiLyQ
/438QEXgGyCeUwtMRGAgvxeeKaCtnf8ndlFNPRusT0S7Roykeb1IJzrFzn5giX9Hu1Ma8klc/a6R
hAsze3C0/wogx4a2sSBQFFkY1ewLcBnLCQ+Gx141Ym8oUoG8shr5ZZYnbZhzi6q2GPcXzQXbX8ap
lQkHlB8ZQquCTZyNicwjxEb49DR2BF3bqtkrYI/5KkgVR+ZCCKQOZj/O18Rj6MNHe1XVxyFRy02z
QSAHRmu2arTBkPnJ3B5Q98eTAyGbzswLPs13hmxg7eYWbV025qsAac1pur970vryH6InfeUOXU90
tWGZAnDXR1MucBaBq3+B2un0qJytoAp6ABjiJlq58M6dmjQ2DS38KTtO8MSMm7GnFMxgJ+KrXh6l
+M0QrGVlfnC4Pdtz/Zi6xmY6PsTxiA/32uRVRxQt+LS2ZJHRgGjhGDMJ4tbI34ttgXTRS4ap7Gw2
24y7tddzEF7CGlLdRr014l5z2ambDwiuzQY50IfzZCmEogO6cxcxVG2hSveEfJxd7lS/bcnHNr8I
K4BvBUvFpedhLlG8AmC1DHeeD6lAZiuE+MbB37TmYERaRT1G8TAoL2XUFP0vnR8plE0n3U4KXG+w
VZoJvVNhGW4Ymg25kn7qNcmr43Ym2YyQBEZZ1UgLrGIG08HaHo6S+lDOMK7Qrpo/vlg4rFbDSOp1
xCworXZqYEh63ghR/jHXV2GHSZ5ZBs8oVNlnNpaooT8iWk75pvzMl0NQ+vx9Aw3TsHOm2vgdYpEb
bguzAxmb+FEEu12jJKLotGgQ4ABIguL275beKjj/7JkdunN6/kh3HL+6nVVww94JfYtMnLK7xrRW
O3OJOXKFaF1qsAp7Fo7yMSGUrzl97rXN3ISLGLiLbUhmOqA2yBjoI/llw+VcJuOKJ3cq44+npmVI
XVer6LnCDE+apUNMQZ5LHWomZR2kMrwfizZqf6SKTyi5dkXom/WVJ/Uc+BpGLDqO9RZuG/9hq6aw
zjumVonKIY3Zg4stl4CqkWhwX+eLBFNWxPHlubKTgb0/vdEN6FhQFP37eiXY7g8RUlD43nMwtj50
sDPDUpXLnSG9j+9x9LpwlXGGsdgBTssoj/ucslmBeDBg2N2l8r/4i2nVO8Xbwm6tRD5hAlKZPu2H
TWTcsSKS1dNnHkt6CDHNC+auq7YLEU3QD6Zp4nfLrEYJuq/0aazKYhrKA1Zn8QqWpbwRDI8Ixari
A7FVuq1OCk0jFw/JrT7zsF55UNQHz4KBv4LbGW1t1zhcND27N33tYNGqJ1BLPJzwwSj3C+lzX7gq
nU3y4V+0blFJB+kPKEXNrQ2FciYqB8dH10GPODs0xjT+muMSSu68Rb6bBiEnAR9oD+/bikfxAONO
RI8JnpK0VV2m3DKl5og2apEPOxWSfO1aVf+rMRfoLkc8ufrWJmaKU0mqeFSGLsREqjyp5OPbzsUJ
uhzazAud4PCS7yNp2q4pGBNfGIc6PgQZ3pcD4N5qVvKxa86a21WQR7t37yQCMNhhnQgmj8RjpKHd
kDg2FfxL5yos9TqHmUlYydoFp74WRWHIIYO/vns+4pbacHBPY+dqLmTLv/JOfZ9Uf46obf0pxuSH
j3DBi3s5D7u0Bd0pFsbKhXUMbJZwH24NRKRicJ4ca0jjgLzw88smnmI1Uf1xVouawcCAtETFkkek
unAdDmLLq3r9dHvC6LmtVHrLBSeyAPCTZAHS6hD5fTxSbytuOqbe9H28zKv495luWeFx8eck1i1O
L1zkjVxHn7fC/UklxVaKoGY0TX6YEiT1x6p0RKLM9UnqB0ScApK2fTKsHTeJEtHeFXF216Qq7SAX
hu2qB4/zNppvDZwQUOZ/Z/0ShkjAHWo+klzFDw32OxhNEt0U9pjvNZjdv/kOE5Pw6wuKcJg0E6ow
LIDw2q79wseYDB6AxkudiSUzCnn7KAzFuupUOYyBFd+BjkGGimcVbTlr7ChGNyfQCnEJY0KjFD8l
uBwT/EdEX2Lq2jhQ83SAOICkjKwkY8JMhPhi0ep8syI8wlJF8+pbsJK9c0s48hSU+F7J8Q27+Rj9
xPIS15sT8rW9zUfxRl/blnfPyBitS2Lfp5ustC6FovTCnBHU8j4PTOvNeOI5sjVHyFjEKG0hF1gB
4nNiZxo0JliqN37+PHMsAEMiWJSH7DqpbAdSkb3XvVVrcrR8eF2eOVihn06qi3qa7TbODBOJQs6p
Eu6WL2DwbgWFLstEJrNM/OwfEyKIuOtPo0OBLuAPCsSLl0FO+nor+i99fn9hn4pgc0m8lrqpMKf1
mx3d/3xMbVtFFMwkkFSj3FtxO80yU0OsfbbB9aRYRVM0slrkDX/QW1aYZ5UE9bWrNnIPskqmMVT6
J9zmZMTCCkckuKhvafsUmllgNPuyGVO2+pR6l2Xuq+lkTxNSLCA9v7hNCr/WrDXdCJxH+mH2i/ks
nBYwAmUueS7ur4oW8ktJmy3a1T68deKv+0AxWGw71mDR8DVERAScb/OFC1Q6mLdldzhsilXWQP8D
O0/GbkdmAm76EWCweEw6GL0tdTtnvXwmAKNJJO3nJGjMvLSf993ujEo9h3LP6+UObNP7rAQKgJn/
CXZYutCm3/65p9dnXHEwCK+TptLbmGNtX7SJasNsrEA0rsuI6CpMnlVGgoNoC4yBhjIuVd3snta8
WOcW5nErqx2NwRmA+V4pl+8hBYCJ228n38kFT8A74re+9n9s5dL9F95e+h8R7c9/PsEGOMv5AyR3
0epMax996oAnXxkDlVm4uXq1PLJYKTtpVfYJw0oq8kiKNgLwx0L3QD9sPrPpCcFIFl+hTZ2sULOl
t8rKUwEDEiN1BiA8EVzJfXP/1ivzdV5M7Z99kMHG9VhrmR2eXCIyhm5vXVGsYspS1ccnc8EK8+CX
WcDIIUk+0mGM8h3Wn8WmHI8QTwl8pGbYc1GG+ShYLZAPpLBs7OtkQGFpMqGSmgnanxaCeBnJ2v4Q
UHnwDymYmjBwKMgt/yjlebbnbIdQQihoXTCUFomZ46DpXuwltsYMObtY/C/z54981NYJrQX84rEJ
ioexeI+N8xEfhaywx4SRkNY60VYnlhiiEe2YebRBRGcsc/xTUoSOB83h0hCfL7ScSLbvIjH5WQbx
Z4vhUmux1WvuhLneM6zZkhWG6r/t/7tOJU3C0WcxWktDODqLBjSJuHk7twoZpr+s6TpSqxcXCUy7
V/QXDLvv+Jiv/9JxOMhQpuAx+Fajy4+LbKa2xT1J6imQ9wnYTt1bhEj+vZhSWLj9kLyb0OdHWt7p
i+apeTmMb/vgvBDt3xTZRT496/nteXAZjoyLJEoduP71DWFZ1a8oHHJ0aSiLU4UyoZqJXttKKBln
sklD2xw6YdP/nUByY8IF/nT+W044TB4GOw5w0DVr7eFq3wYcpklWzGdzizeMx+zc5fyJ7k/pK0UX
feF1chEkjMFs63btyItbq6G4yVw6KJkb9XpmaSOiSWxexFeSr43rI/MjhV/uquQ/g5xaXRUUhKIB
VYbeiLB0VLw38mlGews4+Oz8xJVsbgfd3GxwU8E7vy5QYthgdtswQx/JP9CljHjHp7HCfrVQYV9W
91nms/Jov40DhvF2ar3twKBRjs6t+hnqy/5D9qUGVZ/xxD9mmYVaZgTf9EOkec8ve/f+ijCsmDFy
7t7tGVyXk3XLtlY/XO87ak57k9jPjbvE1jEAfLEDAtx+vO/XA/8mwVQ+gzGMjR8uNTXV1uRuDptS
PfZOJSeqBq10gv8tp5zCyRy9IhGDSOzRzq2v0VC5NKC6DnQNbrQxb7VMe30qHWJUaymTGDbsTxPP
BZcRBd2z8dPFBMiUaUhUuisd07aat2zJh85Nby0XIFmc0kY2X43K1qxkb4vWb3c9dmKAyW4kDIm4
ZDQ+LKnwLtuHa7ygeExutH5MFiOPx87RlvDJRM9DvrC6ZBL8aXgqCfcPT21QLl3Bhn4nvpO+tCBA
kTH5+g3/fSqKkWLq72ut58Plmw0uSo25I17crJXqxDUGRBTxJXsb+gZK3m00Z3LGxirWQsQ0P5KF
d14430/T/KdpfUIiu8pGrQ/pWIguDjl0LyV3XIvbskgWq07ETXCPaJjTrNvHfm0atd2NBZOe33nr
YI4OcF9mKrC5uRjcBXIR+xA4xGNcJ+N74eVJvLeFWWk7jOqE8eSNv8LtdlLP6cP/hoQLR3+BhWiF
u5BAJ4nD7tHk/u4B5eAXQBr9bvkBytk5dQkYpRgFLPWcERAsucPu+M6OMocJIszVuHCRhbY0MN6Y
TReaCC7Q+v6ePC2ttphOpfuANAXHMJgbrW6LID4OYKXr7eHgV+YfZauIYMkuFlAFqNL7bnpYbs9P
w5TVNeduiFoyOEsrenjjTZXCCjP+qVG03dlyLdhLgU79UsYr9pH4WxKcWJasUg9239sPJp7ZKJSY
Vei3MxhZzLlO4N3oCp0t3McZ0GiXqDtlGRF83JkFg3PnCgV+UGK30jvIwl7kvIgogxNyCE/789jS
8Dc0UIwKmsPTPzGpRJfN4JKvHiaD/NvrkuPvzT7j8AKIpnvo4CjWuEiRE0cOlp2/Mh+lj9BmzHlx
2S+xOeXegLV4c55BNcLNgfa9mRSuO0As1sD2ctN/9fwI9iZH4R7V3KAxvgZqLP8BqNFl5dAl6GhQ
/1fj8jzuvQoPc4wbVGy6dv/h/GNddzT63ZOf0dfTOIMVudecnoDbxJsm+zMSS6r5F58Agzr+s+/o
9UzyiIlalKEl7MRD8ZAgrwEq6tyKqVC2PCucViErPItZncIsg03Myl+wSSkMts6KGd7dXHCYvLVF
4tPZuT7hzxVTJ3pvFlcURYhQBrK+w+9PBJAAbKQeXRCvjYS7MWYy/AWit/4qGxyztrpTWNqv4+ea
joIhg5HtWgEwkVNYNdsWnKQltpfICiTs17WgYlAviki9sVXMg0yKuZwBZfvjYn63jihOPDoU7R4F
rVjy+5oNzL4qQNyvvhVzfSSuXkG5RV71URmazXXTCKJDMaFF9glFzfqr8U8K7O1qLXx0E2v57a8d
kvPrKaqhujrXKASsDLePJtop9u37GJqAicPWdvJ+zXm8INE8pQzcnZo2cdlkCNWY/iKuzzkSeD2M
m/PsjExJu2bfOs+RxDUI5Q5jag9Pr4DTIPv9nIE616OCunUaLZxkT1K7Yd/37mmreawW90Ty974f
X+EvxFJ5Fb39GjH2qb+OO8CbWmb7DP2Y8Y8zl7fdRAaSnc+YRtYd+nFTl26nt/7afJb94jCdT+at
GHAEKQHsOcakW3cO7PUdQuYfW/208m30voCbMCCpysBxNtZg89RsK6sYgPwt1m4IGjWa+BxAHjdp
zDUnh8u0f8EMU6lNudNoXNJptpvJbjl67L4XGk2WTPxBauhmZnsU4M65AaYbDJQj3xvMEYOCbPEo
nTLiicK2rMoke7p6XV8FcjW0TLJaAEA8qTeoKC2k5zic+SJ+9KJ6B9ZA9d858OvfZhkc3KbYJux3
cXJBKOdonMOIHEcQtNNRBlhpbZplVSOu0DeprvLcu6y2xuk6vVBSHW9WCYp/2ToKhMdVYaBfkiEi
+qj1Y0Wj0VssoHPLrqbw0oh+E4t/0tQKR4M3r7eYp3B3CUPN25qngmjpv989I8u3shSfquwPqACw
EiUBw1pQpOBBisnJpi0UTzcXis/YpidZLWgj7cXblrkpg/9a2cPOW62G2uhSUd1JgklzrjRW/YZE
RrTetqHxAycWvo5OQVuVj9Ktq6kx+fgTv7HleIZmhJtqHxpYLr2wNWePVk7OXnJiZkMNZQhlh8TB
Ck53k3Eahs4Cr5jy0BQSLGjPaFaN1GMkBCFPJ8iOtQFLcqHpiVUNomxTuvvORp47NI+6WWBKYKy/
9ZIL54JQxhI37tnyorjYPSj+gNj0OXCKmk5+p/Pjo59y1yb/xcAmGdt8NtPMOFWWJoLdYJMj9eRa
JJdg5boTGqAPLDuwggZTvtrMH6cu9i5cS2zeBBLtevhqpIVzezVSSNLAqFmX0TDyznk9j86ceklt
uRO1TEhxvB79YvUxPImFnZbdhGnMA9foiAAMVH8evHGpcOY6Nf9UQPLqhuKJ2XS/bylvu35N+YjF
4lOcibKHZGgdX98n9UHruIsSdt9HKQXLvfVH2UYoRA40S2lHiMKBkn1xWT1IXTz1DWPfiVpmw2KG
XwzgL/WOIgkmf410hoFtReHyuRSr/O6YaNHcG/BEPP30pRtEF6WXC+nlXaWvRuxdLCJ88UtrGoow
t3lH/l9c/qDpkad0oOENbAVTgDBRDwZsDvVDL0M21DUafQoIRGEeM1Le53Wn/isKJsvT5O8X1JA3
aDNDoJCOFvhIIF7ADW1nY6ZSZIwceOqbhHswJ1QFprcCYR91jVbX9V9Y51SK/HX5WNlmbulNioeY
wkmFH3GkF7Ual8PQMzhy0m3EyhFPSgHi5Xd7iPImVGOJxpJEiuN5Hljov6uzo+DTUc51xV1U6uLk
Ncj38hFMRjT6vhcFrZXmw70qlI0/uVC7cFyr/WlCHXs1Cq3P8pKD6VlKbbeknj8eCOUT/oSudUr9
vf+WqE1XezGY8yHiqH1kZO9iduAvGBH35PnpN4lEAMLLmD4ruMsa+HLqfip6jJa2kU0x/5DgTqbr
qJoVbctXYHv98E1rbkmvliem6SZbSzvdLnAOGZBozijgcItTGZKgf7GFOaHAH3wM02Voj4EhLYch
IR5XEwEUuYzrPkPt0XdMtmScT9J9NPUOKv4r3pwYVWpkHWUie1ErA20QU4sub6IzGLDpJoKkJkX2
RBRgiEia91f+qsZzn0yyfHoE6kqETLBXWdc+H5+Op+G2y3Im3zecv87QWK4CFz/82t43rxCZhmef
agc+XyMYJpBjjwxIbCPQHs5/GviRGcuRlexG04QFwEQ1Y+hqVFwlES2wEiQ6BEwteTVMGhl5rVs/
ZSB1jjzEMGPMJrjWIaRkafp/lrVfRb4Df/ADEnKF7HzMJkFvHg/BmTt43eACd0NvBHjtQ3OVkYCz
0dTE6LF9AIJ8K5YhQnwj0CJTW1Ohvu0tCxCvgpBJl8ICyaotF2hyPe0h7N7lvLWpfCCY76xRTsst
LYsd8pKqmFF+40IpRla14pg7s9+AaKgSKdF9oMJPPNN2Y4craKYlNOx9pYDeuQqYOFGv2BElMVhZ
fIPTGl065W/WbcHRelXrFr1PKQL+0cRjhFiBvvPlRpOj8yuOrjQiuHIXVQlZ3R3EyrkQNcvznWRd
7OvH8WUmTS4NKWFv4roEp225UtHCsmbYQy/f0ZZg7G3IbYXR07AvWaoBPYDyyc7/c4Zy9WnZgmYs
qo6PZzfluAlN/ILN0p6RVfWiG27BeOnl2Oh4/v5vbEzTahgQaJ9pptdZYioQ8sIW0jsMvEmMVj0n
gtIXQhw2vpvaliBlGF63Dc1ORU5NES1aoa7fB1yOXlFXrvhLsMZ5keAuQlD0PIG8XNgoRznzFaoe
RgPCaOOw/tQwGo3FrABXLc5/rqkIqPPc3JpYfD4ObejrFqhKie+m5FJ+WXZSKphkSDxDdPmDKbNg
iudIRXEk7LCc6jmtpYxmLOAZ9VMNGWLwV60yYZLGQW1FlYXP8D1Zkv7OFQ04eP6v7GZbJPpreZ1v
ZsJQf9+xM0Wa9DZ8U2Pe7mmiNBSsWNXihgz3mGBi7g2EoKZlRFu994CYLS3yTl57HaOWtRJrvCwO
J4GryKvFhs85U1Y8WFchC52aIbkgdaQAErjf3LIsk01aiegZRwfRNlGGkXbiJAluTEWClm11wB95
ybiR39L4o3qbcKRhELLAnIUELhWEyePurIJcb84mUw7l0+IvsvUw0Oto8Cf0KuuS2CukqyK+HcIM
jPnPBZjV70pdUv0g1I5T42amgZIbr0yKA5pkUw9ry3gxHXe9GmTlsr0oPleRcFm3gsMKXS/PY1ac
+hTwxM+s6g6VbSVNxM61bgPwwmZvda84IfOin0vhAQYvhU9jFz4PWhPNaxfK5OdS3yTCO7ZldIwA
+2ybygpEyVuLMdDjFWNN6L7OIkhyV3SBGfV+6LEe+GoLwWdNvH4FnPwZpglFPu43KUFn/O7/wG5X
s6uDg8rB2YDA/owhq7aZ//enLIMMUuTityJdWpVEKTIgFPa/Dwk/RusfmBvJh2FLpdHcOZ8pYtyv
SjKW1fVp2UV5HjhcVFiYsk+/OtAe3j/Q6mlL/kmUJ/DrlzkiOxzscvJGCSR8T79/WWzjosVZ2TKJ
L5kK5bmOXzvUO9WjtbZxG5l/KDF14pwRdfFi9JYr0C9mH9qqy0kiPKAoXvLR7Tr3be1/qrkQ80du
xnXNGYP0hJWLISjUy5+RxV2c64kr3jrl6ql/1X6MOg1KRmbZN93agEgXFrJSWoNxA33ZvdoTP24A
kQQQTuQSmilIjC3KuQRGHkPn/udsD885k9rat/ZtKECDJiR8Sp7jXSwXwyWXwdHcmMZ3DOOTw67Y
hR9zB0cQu2DKgDG9/JQgRM8A7EzVolmebDd7ngBzQpp3Q6k84LYpaaaQh3h6ICz87oArtmcsoZ4l
BBqozjOOhBkIO9HUY5y66IhywesN6U+sX/6fSQnXh4BZUnkLfAJfUJrAC9CneIivpt25m2BkBsx4
nx0RT51vynrHAFzqHWuBafFEBnvjNUXVnkUvIZOxO07eONUbGfPgCix/ypsGQS/9ohLeo/0ScTAo
QQurIySqGHAdngv/OxlVqtd1s8ZsZ/7k/3rvlRpubtMncN4S37NgPJChfAl44D3hhWDgAzHjADNS
5MbU8E5TBOZo4vDyIScY9BsVgjZLQcNSMpjcnrH3ZdGH1Zcy1EXz9eFvZ1aetZuXZX16bvr3Wrrx
/QY09xKur1t2MxrH5feW8mEQM9/qHxBgu71q06dZHS08UAxnSJIAPfofyDlf4iPLi3l8ubeg5d5d
+UWzo+eQc0qg1rPwNfQ5t1src6+XSgzK70/px5wEn/yYkowfsm50HLPLWFzgdh8Qpr0TtA2SK2rs
NnOQyYD01YiNRKjJwfbeq1x/4r9GV10qoXnCDjr082+mR6tM0qKtIzHbuM2kK29pRkGxPpCAAKix
0UhhUXMuXAvBGLnGoLlW0KB3ZKchwFqQCtDQ2YegO1X5nNEGjTUoPUQAx3DVfexezNGAvJQgCEHb
nvQsccWxskMY4ldbat9gKTOaInaNWbUPpr+sM4aSr+ghK0g38GX8lIZAJyrl/CpwEHxqoN/0QSbd
cPZwF8OmIsO/P7u9IsGECPcmaBJ2bZW7wDbAXsEF6sehnPLnMtfxw/AhfWvfv0WV+P1AkF9i6W39
rgpMZFPCTzHGBwFzQJQ0yzKKLr2sG23gxMPsRfp6MYZZN2rUbZorERsNtGb/eYiikMeiwQQZm7ca
MuuVt2h9BgBoxADZem1/SRH6nZAeZ+a+/Ri9QMEx8v6XsNoeSp3g2/wxzzSHoCOQwL/XxvH5uvoz
KV2JypvLTBqQamg8aehmIk8j5EZNYxY+5dxs6GgU9k+LaFYY/Bfsh7gSp+Qt2WpoH8pCAyO6jvAf
cQQRx2qq1mxWMkrhDDEeyo4iNK0XQm1Tc2IygY/vnW0AOg5uWTjnoECrngYtmXW1IlZVSZScKYhB
rxyBbRV3kTwIpEXqJpsmd4+slHYL3+I7WraOifnDxAhUeEqryJUGtF+d7YxQsV5UvWLbk89JYT/5
Dj40LqkaaAu1jqB2vEVwr0RUoc5CgIBEe1h0kv55tu/B4li0G3abX2897ZN28AFr6mqoskr/dMOq
HDkc9tAaTYt6SbuKZor1hYkFphKm0TsFWe1ZR62scLA55Di3CFuCIEV9IelKxPiLc2y5EJZa5cj0
gHdy+qRgI6YyngmnXsAJmxOaeWC4DROdEliasRN75nR5Emr8waCfMlOFn+uME/que2usEdfW2Lgi
NDxJs7Is/nmuhMqpNzMNOW+IVp1j5qBplQXHnc23I3M+TWRYPF3lDtjHn5mH3CvuKuaC+J/0Yf/W
PhBl43G+q1LSdiln0E/g8e6Qm+Pf5y7/82tvG4tTVJm4YpLFpCD6EibSae1AD7KvbPg5s13Oaory
4+yQWLAckMkFQJbx+oFc/yg/oCDY8jhMToJ2vx1q5YxcsP8DkI4kwKxEH5gVjCo0c/3OCdwsg71K
IQ0aaob9h241uDoN7TY2bkUD1x4Ixd/lcmh1+yjo/gTrYPuzLKjkYu1P+Tf+nY5Sgmww5MQzyyF/
eTARiqzSznLYRYZpQ8k2a1QFRiZcp3GahIf9sEpF+TCj1j+kTUDa2g3QW5ss5FOrJQd0bMs7XkLg
H7LEIsvlbNktdrhJYbm7lLQGh+PyZcIG8JaZlryB7XU5BOIO73CJdmTdKt3riEFm+3vBOAj0Wabl
kxXkon76dia3qxk3DHVehzjwj4sD+0b+lL5PMBw/cX7sjMZnmS9zEn8c387DX8NY71aoDfOSbTs0
Q85Pg1b7qtbuDAxT32rnrsi27XngQyRtpHTnwnjkK0YIX5n/0+5DbDWif2/0soTxhBGZ52VuPuz4
3oqDIRMw2ReAt3OHs+5Pe86hm6PdvGom9GlKVarYpQx8YOdCAvBZX4SGBLD186ZgcNIBmmBFGEu2
KHDr5B3vNP2Nk4y5xqvOq9GrPNePG02pdKwqivVFtwhFHhl5/OTjN+2yGr7eihXKRLKiVLiWWQs3
1OuGV+7Vyzm3v0kYFspKCi50tKuX9FmAprB86vKhTGfPgH0pZSppMcodd7mNvG2CVC8HYk2FUmFo
tNjVOL2FSpI4PHMBYh52S+2E0dGL5ExTBtplgcFTQLfXf8hKeybGpnetatXHFlXxcDlRbgSpcZZ8
wOpOfVFCwTDErNS9z/iFZZpNpybnCj43C0ICaIYoBCKhpEJH7DEHAf4U+LXpCcprwWP1MUKb3cQi
q50b5xg1ug6ASv3k0NHImj6mGW+8AOb6cTHBgR2E2IegyTkh0Dvo+zJe7j4RauOG8PNMK2CHp6zl
Scx6K4w+zPXL35lWv2h2r4UDO1qs3ml1+lqs0eEkdHq0m9Bk/qdmPTLlSmU+hfk+S4SJgMmS71Qp
ltfgnLfcOkvBFUJ6gOXu6493wSykkchJDxpgDyt2GpBGFnDBI7tFIH6Xb34liBhQ7aV65CHir8Tw
A63lu+YgHyi0GV0TSBxMo8jrPSY7seTz0g0l26/O0PkyZXEZalhNYf7PL3Xa/sXEnEr+XLlilnj3
rg/flHe+hW6lCraCZBFxZ15kZVo7uCWPemLQI7VRH40AmWgBJR/rg68EfvDjmO1NhuOviUaCGAbv
UTATjZ6l4II1QAXBmns2x42wyPk7k1/XhYbfXELovWpdN11dzwm7/h6wxXi6/Xe9PU3EdQnrJaex
lMGDuUgUH6eIScT0+2orp8JTURtf0HThGXTHKc2SM8ZQhjEpHUwd5jfZowJnrsEipMvRQSLJuCUM
jGQFf7deXXlzShebjey0fUisk3wix3uURE1o8swchwWhOLk2KxfT1xlRoimXHiIneEDkSk3ejR3w
+aIiwBKrHK3IqzNX/8HNHoQ67SCXvBb5WCmTa9K0ISbK/SeOodUPDBxdkH4PsbiaJKUbtFU2Sk9u
TEO+mMGX1/OCxfWWbM75TC6MwNEx+TY2OIC/AvdE3SubvZU76ZEfDCbEgZP6Ft3R+vxktbAaF8WL
XtOALmx7UojFlGfDY2qUOIel0FQB4KqG9iXs1U7DYP9hvXw/nfxDlxQbzyxEqZRKr/9Z7SGgYLzV
cE42a1fU8Bjj2yIX1S4B/9d9b3MwtrtvsHBvb7pTZkfKsukZsK9vQLjaKerMYpzV7mHUDoqNS8HR
YDfv6LsSAvymYQmnf6LGkJIDiwAuweqLSSycfoTDt/wyZWI3MGGBJZBi8PNp27tGZLnBDO7YvHL9
oxNiIy6gKz41ibA/SFDuzphf7WxOsIkv8lwZsf57DQqbPuzCzjJPvxQJJAeUXCjqxg8TxjoAAlQB
ULd0fxuVp3lmbGCqCDqgL9lgu31LreeSMuwoVmAnx7WMRnM+3O1y5VownETxCPgiChxMso9GO9/u
fe3iyiQ2W5ZlIH8cBd8/M7ugzaUIG555D+U8+SE7oxe/GH1xvnQ480vCjM5rooRlQO5bgIy6cazg
uOtv8tvj+/RUWtfMfxdc43DStZxNyn6XV5m3ouhTYq2rkX/kxcwqJd2QWrqG/Zb4avFEWJh0Gqu0
vY16Fd8w8vR0mgoTGsQ9Py1HRwR7mQx1tYNbyZ8vZuhRo0my3KTV+vKevH3HBMEzWszrk4KooNVW
kKQeuubNbs5q+BmBof5KqB8RZUy1U6Pm7JpLa22Ikk15PTzptuAAcdubzU0BtV3Ib2y2EnHEFijU
4pwKdmPQx4ovRETSHwjx2mOINJBowWTI9fugF9nYvYJOfv91HiHF0rWAlEFFPSVtDR7qvQT+XUYh
NHXh3pbi9OoGdDWJidwQkCJ0gUm1ZGeWITo0RHXoP7NIlOPZa0KKaWllaTDFnkPSg3V3NWg0Ep7t
SmNyuzx+9yqymej/fSpv9AVjta3KVamNqPTITwYom+whVXKxGpRM4HDdlGkcO19XQwzNIMsoFO3u
9mSAv1iuszq7/xITGGQ8ikvTVz5G85U2SMue/YwUaOUe131MTB1Q0Tbr7K+x5qTD38MCkSDas5YO
taep7tJIiNqZA+cG5FlJI4lTjPOBL4YcppnFNJM/4gDyn16PGQSXuko1Y5uS56ysrbJi7s9JD3D6
B3N/Q1x3SvLjjt0ld+NdWiFL57wBb3usKmbaeTwXtL17d6pb4Jdf9GkSpwmtXrTaN9kXpBtVnCqb
CNm454LKWKAtgG0ZtxjH1Mvt1dsqATMRUwZUbAyi98E73SVXF+Pbv+cCLyKfk7ezATVQftOZVZ6x
cip/DciMooEGCwGmVNrWCMELXGPB/kHtAhm4ENEROCUDbe4Jh8E4WVBjo/9vqQFDJVAV+SsFWkXx
PwTz5hTwhzi1u6XF9/LZNBSOdqe5AWVhaLx9wavb5kPOibTRAHJ2OFUlbm41fayABz5AWzHOVd1T
nUpLj4QEKhjDyd5Pn9t8qqLb8YtF37GEX/4ZXrBeK4o4Y37w6gLenLyit8pIPJ5VKRniBKP4f7Mp
cbKwEmB3T0D17goZsrDukgt7yiSyS7GEv1FnXsP4xb8VQnT1Huaod7js2dWZOMmtG5Nk4LTQSAmf
WBPDbV6OU46K1TSJouisRC4hg6wHj+gGAY5SfQBwM+EXOt+ZPEfCzsHcQW6iexbBUFBX3PJSb27c
5XjX+CKmOYlvZSMEiszCsM282BCi4tCJh3680WATku6CfYqnN0Nt57LpFckQp854bvLPV3oiXUBP
+ia8RcTlFBE285tRiD29R2qi3HpmuzeYpGDphhQLNTa/eAWq6HcdgXE+bEHPfnuy1MYslUybW3yP
SvfFa3js69x5yIY8MmYl1KfULiBaaNMIQV9JDD486qnnK097LivrePz9MkeLrYwzk0o6ytppMF1q
uxalRfAQItIxs7eO9QxrgxYgDoKhmDotU76ZGZzCJhhtpsQw4VmxJZflT5DeV2I3EGL4lNHOwBLP
bmIZvDp7iWQtZW3I7m9tznfOVdFRIcgv4IsoAT7BZ4ZVRUS7fii6u687v6+OlHJ59vcWw25PGU+F
46/DrnC3+6F8J1kL8JIxGXsdBaSQ3R+9+c6n1bJCK+VqqBp/CU+/V9Ux75fk7O78nNW84G6IsEgA
anWIAok6ZAAJOoytohcNvvH5csjU0bkKjFa1Dbc0xq9CniokbNUtZiTWHIPMS9qGFTUXEqt3+pRJ
Nh+YTSW2ewKTT6fu4tHDqZFByTRhveZP7vegri3809BWIXJ2s8hk7XBqOdKUWePN8YXBzH2bh2l5
p0EzkreQNd6Xe0b5og+asrTmHeDFLJ7w3wRF80Z2kixQvX75sY+tXsU8DO0BiiY1I0XnnvdOuXF9
LLR3kvGoNcYvtKDio+F73Qf7AjOnDNs9cnERRXLUSIx4ym1vXAVchjhrj6fg/De6O4ZRSy/pUOe8
nkcIOA==
`protect end_protected
