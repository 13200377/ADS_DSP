-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
LjD5FWQWvP92K1OsSuIXAsp4f3gZHMrNGD9DWn5HM4E7WPYkNIYImppvFXJxAfAfioQEkg6Xs0Mx
cNRpB4VTyDnBXUYNfaqmLZtEZ66s7anQRJUAuwe9+0xXbNpbO+1bjozL8XOpu4CWeVh3XRQgKLon
JRnJRwVWX5Iq0sWXmREGCvR+n39W5hzYe1mdT3a3iVaNNfI/PaX+N6SIm5sXe3gC8iUJkUQEWVAs
UeHay12Agfn6CvJnsLa/ipffDQAKoCRoapolZsU8E7ZYn9rSVzXTYUWBYGZ47vIJmOhMxI686eux
p2njlZc3BiesZ5+IoNugxaC449tm8hZb7IZ2Gg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4288)
`protect data_block
vH3BEPfYoZA+2Uv9RfdI/VwM99PJiKNOfpyx7mmTQZWxEVkJ4uvoZjddJ8YChKd1h0NG9MOmJSha
ksYHBhBfYWtzgTHUEFuRAJo0ysrHDmNQg+UTAJ6u98StbQqeGdFOj8LcMCFOXvLOSkClQOD9FB6k
9cn8pg29xu7RM95AwbQXKVtj0WMpN6Y09MHy+AAIZyS5NmJNPYHzPLBNNjWrfyJecBNxgbhzPaI3
7K9SnE4yYIwaLvZo0clRJl8f7jmztLlZo04tGmAHcSZ1lbbuITWxxfrHZV6xT6IwNOvhBVHc7ywo
LJFNjwsOgMAgZAXFmhpzgbwAnne8IBOphRv80cZEIOT5DwHUXUWkfeAANhQ7Sepm5lvnBRm1FfoM
Vd4VNfF7uilMAyXRP3THb7f3XMeB8Qrofx44a1eYVu2vSOFJ2YjND9CZQ7OirqqPm6PBLhD5jPO6
KFF6WuPGWsVxj62tOE3o2BBpn6Cy0Rxg2t7onAAOBGA0T5Sc3mHhM4oaD/k3vd0rEhcELTOaaNiC
R+ZOTZZ1q+45n9JlAy0Y3HpMkncurc8xN1CToY+clT59h7rAyQfLdhNFrmldQtBEMAVyOmJ5KqXr
2zJHAKXrnteettXwshTRUdEvt5QL5p0DJEjevpryFH+NUmmMnifsXs60VyIaSUr/wcxwfuGv18sw
MzSIiwf8I5856u0RT0fbT2fYT25teymUMgrz8arlcJkxfwPvhM1sodUjl4tAnMue37GxEYQ4VzvH
VOHulg0d7bM3Xtt0IddhN1tIvGTUZXzyGRpDrQ2p1Kdp3Ooz4/NW2sVd08ZhTpcwC5fVsllH/LYO
atXH/Un3oHELi+F5D+h/FKs46H4++VLGr0RSW6CwqOjoKPPxrLQ1v1u3mQvUU+eJrccQUdx1nkcp
eRHEv5am/EnPZpqi6HZlLh2kjZFHByEGAKRz83tgl9J4EZUfjR9xgUIW0fboRaJVF3l4vOC5ULOh
UMVDAWawrat+JCMxc/6fcfJbk8QujgRBQOUfy55T6ZKg1+Q0o7lyA+QMsSV4HS3tCxw0CpLZn1Jr
yIBBJrnOLYudukFcFWCX9GZxLQeTDqBEQe2wzB9fWzb+QcLJeBLZsd07lS9/U3ST7D0x10UZXOlh
7gkxjoybAKXTPG4oukWhAtOvXc3e/DTM/bDsz51BpQQWygI0PWLowTCJ7tiRF9zPO98dQEtvFj83
EQ0WrSxyyEqOpTioGKoOAiPORYDDEWeZGq2KptRPIBxT01Dyj6SkABaK1e+Aueqdrzar9tsLhxst
cznuZz59LVV1pfon04wlAd9Fz6QmVjYIWZwsOu/Z3zdD+LQipp+3Wea69c1vW2zrUYLOomj1FgLp
0z8tvFTXWA10z+5jLlKFVgvKOIhjAeV0iLkslJT6EU9kGYmwG79UA0jNTFBgp6YJaRqU/SdzLpV+
7t9Y2uLd1XJhNXxcYaVZ4h+ghgfZTwSRwdc3b0oEGHGdoNRpHPLaLZqgx4SHjwkniKfPHbnJXxOO
6mgIMVNS/+7TvFc9LeS0AUBRZYGeV0LB5szmSN9Rg+8x8vFZsqdK+T7ZocnwRXF1jSznME9/fIR5
oKOnnfD0x0pj+7Sy64Al4KmN/g4AdmAcEugWD29CJm11j5SAuEVCGQKaQmZsxep9gGSibuP/HTkF
oROAtnSQFb4PIP1pGIO06sPhVmi1DdWcq90/cADht2Q/r3ulScW8BiW6WcmQ3L2zbbVrcYDRUC56
gMRws7qv83J02HkdA4/Qwo2hah89A1y2I4IRQ9tv8WwC9fdOJHDiaWKseY2tHTWHGkrAeMwcFGeC
8LwzxN/u6TDU1lCM5Q4kse7pwQxHWCSiIKUN0OaLBWxBvtKak0R2/RlHS26ucI3qZZNnbe6TWmXR
gbjxxnu8btw7y8yNjzwNxlaJazg477DVL724vM0Hc0JaiGhfIpZnShQ2ms8ExRnJUw/fA3kqgNDQ
oTGUm1VVLwD1LxRcsD9xbFq5YeN6m7bPVGixvhDSrHTK3wI48LKLMlHsVfPY82pqPswgMNGZhVex
RyDS9NcrtC+KLYcmBif6V/VLNp+fEvUp6aK63UVRjlKNw5r6wHp7P3nKrJoQO8OfVqIFwPOMIMlk
t19Z9NH7Rganygs1GGiJGeGyW7U7+qxblF4CGVgdXcZ1OyrbW6Z61DnuEDsWK8dfnYvJg2IipRqc
zIP1Q8LZnADAf7P5/EweJREI9PyHN9WDr0c5lD6+0bfnDK5TtnoqdqqW+mnzCbZJer7WLonEtNz+
5juod84JyayhN3IR06O2HRoqull2sRu6/ahB7kw86kzSsR/SiBpj4bvwR225O5pHhYRpshB3r4XH
/LEV/62anzX74JXuBgcRpunqNkLByEz9TLVa2Pp3mDEQaMsFY+7xY/BW3l15Pb4vF6/Ooq1xOHz7
vnucPWRIn+wB7zn0/3+a1ccxpUFObpT3Q4KF+fAKg7EVsAKzpy5/GTxjAFyXWwIBwWksQgooKs3y
Vryxstu87rtNofq8wyS8+6yaMwEI6dd8082Oapi2PomoCIDh74JrrNice10D4KV5OMG7/f62QKi6
nIbzu/tT93MnNKWq26KfmGaQqrTCav19QZsVzKtJbAeDiPYTcl1yf3miyPSzh1/TXeKSJmkvfbFZ
QlYR7ZurOI6zSs8RkDdIRxPA4goIFvnXac1t7eCNQY5n4q6CVd8XxW5SfTDj5Y1xkbf59ZyzL8/3
AkfgErf3tYUWHi26gnf3xCTMvEdo2lZH9W3JMOjkqo+LZgFUgxLxgcrXAWNYNKORtyY/iVj9nnnx
vYH4I79aShaaa8v4wgw4dPICaCg1wlzWI67zfBZhTga6GUxb6ALxnojpn1h9mx1TIJoY1PYWgJU6
iQ+RSmRKudSluWgChaWClGugV77okU5mORiP4DVpmmQt/bsZ+5Ey0pqaIivXIP456tGELBQgbJ1D
jfGQbOV53ILTao4vD0ebB2QvKbvbaBirpkDP9SgPPEaBdFMXmNaGEDRRW3krMmhpmKoYJ9fJSG5t
kJwSNRiIWvyunj/L5gGRnAoD6ZaP2h32I/3s5jxEGeF/UlAkxt7FbXfBO9mzulBZAOGKBcv8YbBe
Iw3Z5Bm+PrqXQHVwgjBg9WKyaCrte75aEW/OPFzKG3NpegHoQkBbv8RiLF38uhQkjk1d74CidSDw
w2ZeOCBDDdoQNvyC57TCvwAEHPm3PbziP8ki/NmZ7zhfHXXHEO9OFT/v53I2OWpiNJhTzxuVF4vU
CDVRpiH+DZs0xdIfOJuL6kRr3jJ4I6pUvIjs/qVzybiHpwmIuJZfdkXhg38ex7511l5123J+6CRw
4/cxitGn2Q4jn67nRlTDOtXh7Q2WVy5umZlfB9FAzEv8muemKGoEJmrIBsj/sJBtTgYG4/Boiv57
/R64BEGN6b/XqBDv3NSWL7I3MiehuEM5sB4OhJg3qwjTV2Yf1XuHVTxfUzXapI1rhfhVublqQ7HR
+kCRoPWZt9vvIxmnZ3PZiWCVZ5+of0DQ8lXVYlY931Mf+sFhpvaNxmCh3xAFfAm2Y8OZgZ7r1ood
CuaZ2VU4c6Wu8oXTE4hEymDUq8z42a1PwI27PlmbxKjFpUvMgvLPDWaX/Gl/vlWH9EUtZviINeef
/ot3AxHXa/sYhfsbBBNw+uromgQrPPKUER3C8xa5cwl9W5FzYMVIkSQT6e4V+ku658aZYC24FsY9
ZL8QLsFQ/Utz5xIa/0pGyQEyE9/s8VCBkPtm/6/CsFO6zJ/OIFSnR5HpfBi5UX6DVuV/YCqBvnem
RAAO3M92YoLve6pFnLH8rsophWkfDSZBQRbwPkGC4judRLuUgO/7S4MYkDN2gdYIzbVzBy9f8l0T
LRjwGFNhcnEAsJ7KdStjlLrVF0OszmHkN2ibb2UXFs+/PFWTmbAJ+CMMUsnO15VPc3Pgdw0Eal2I
ob+0T6Ui09emEavf0qNK5MTm8pRVcvCsEIqweGvCiuJaQSgu3Xj69oD0rplWG0i0VapwfRcoWyRH
ACvCD3YsXIbAxGOg2sQ6XAUdPc0VlTQni60zcjQdTNgQw5veQCdzXHm3Tutl2Zm6pD3vmnD9Tm3Z
c3QHbHB/+33Ju44r7UoK1j0deavSfYpQfikVoIF/cgG8gLmSGkc96DphwSziSiR2ErDHJHDaCfBF
on3A/nFPRaJDWrNHmKSuqadFhzxKmG7JQeepAdWxDWJgEkq4pdy3HU75Q01ZlA1pglR359GC6YxO
Z+8wNCyMXNVa1WmE4K7ICGUkfDKGF0LoE+D4oA0B+HDzv+SlsPGJ4/54cstAEl/uuwYO4hWYcC5n
PL1kxc/sMStUNmbOsmOIJcJ59X5hmQSeJBvGpc1N5UXXTAdsoy8838z50BHh1eo7ux+zLL96EIjO
p0qKhytw+lZr6ZJoE1SMTypmK97BXMQSukQQStxT0os7wTqTpz8PmcPvzbuvnr7bcGw9qiP88bVb
Jk0dRXMg+pnW2FVZkHSpTxt08kvvtCd7D7/7nXFwoO+ClylOmz3EvuukiYXqJkaJ7RPIyxb+5yVJ
rKpDvc7laBq+qSfdapVxpn0AZHH2Fr6AzVrCt+/hUDjj0yqMfitGMO1oRDtPwZ35m8AQrjGCwCpr
l2LyT9QvEr+8TFSRKkDaOi6gXaEOdLzkSNqyi0xIhYwSAxHuctWfj6UgRKvUm8Fv1dPG1QgTzRB7
ET8M+oO2tI3d2LZyUbKNqpIluxBQ09DRApfyjah6CLP+WtqifbU9CUI3y4ZKf4RqkC/rVy4/V18M
orYJVkRP7vCD5IFj7MY09SuUPyuRwyUOllvF22xvR+PPq59j6YDhF47gShZhTsYOa4DxjtC14k7y
dGnRNf/nuEfb1wh400BqPZPx69YQevIKzAy131ocsQPrAdZWeHcn4UUhWJ+IqtDaJEQUq7lAkWJw
06Q+AXmgeV4hhDPyNKXowckDV88NJtxJb77EG7hXGhzsQ4uz2CbzPdUZIZ+RqC7i19vOMpUdbSmp
ShFSViBA8RH8sOMgGFsPygKZRTy3b81OAR+gkMV4Jft89P2HurrwwBmqj7NBZB3+1VoIomoLNcXT
1ByHDF/VS7rEjWELiOey0joYWOWlsgv1bGDj+wgOhKtbCRtmQq+vk54xL4yTPybgCyvObhjnJbIS
qm57fkmbQIEuO/BbnMiF5Ccc6w8WLLQ9LNraok+STtzy4LlgrlZNtiaNyEIvh0exUfR+ppQwXL2+
Udgu4PYpV+4B0zvFG+Inwl1I1gE6B648e3nQdOavwLxoJG4ssSo3o8Vybnx3pD9o1CcD/JCHLxee
zektr/EQKfgyBVdb1fIgnoHBpj+wkSyRucyPKCokPpn6MobhWYe+WWKjCzcO/woMVepFbxVud7Ob
5mzppOF4T0jbiIHMYxySJxFjUB+Csn/rH9SWoetKRBllq+6HMphj8i08t5OyhnmSqikIOUTqIjY3
Oz1wbz1wKye9vKmNWqahGGrFsAkJEfx3KPti4wLADyjZgIbG5g//Z1AIXBE5VCN8DGJd8hQC6V+e
l1PlAsOxWOtjb9hd3N05Vxp2cuaW/IOvcos24shqHTVf+FTvVgLrHck6BbBoe0Nd/A/absI+E8lD
OpByMIrs2k7Fu4SpY6nhhXLasDu2K1HbCaGyBkt7gs/jvp8ThbxI1lx3gBucZINK6JXI5wMrOFXz
C5iMdvPAedSdoeT66w==
`protect end_protected
