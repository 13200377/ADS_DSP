-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
yCaddbridm1ucjM1u5n8aYlMlQpxBBp1+ROzF5yoPPfEM+p0IZSfu2lH6tB3qAhzzOT0BWI6N/r0
Ba7J6MTarZ9/hiYapPvdabXZQRucRAw7s7uM1oVawLKOD1lk+cANI71RexC87x/VqoOJO7GVtKjf
bjiseEoWDQ7cr52Z04E94zSDvfoTmoQB+R+ckbQB5pcwYvOgDgR5YOq+T5pUYZs9iXwfjBcVqW6d
hxIMMa2sPBayYRlIPBL5U34ZVpbHAqIx1iueGG61P1GbolNlOQreeci97Gib7/MFDgQxtF31TFul
1X+CPY569FK2DnzrhYyqOCsV5AOLW1K+XzPVzA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5744)
`protect data_block
Nk5Loe0jtrP/qkh4Z7ACvPBCrUmKMFM+OxKVyM/DcX1xjlwv654MOTpF5wDBScqMPKB3wD2GJiRg
3NHwWgZ2XFUjfuro9y3b+VszuVTIt20/D4adRkcuTuq9yZ47hSEMYdzAsNvufo8m/xZMa1gJ+GOG
w74JR3zA15Aj8uisWuHVxKMrhTKjIGDvWrD3tczO/Bxvrp4GKBhShou/9ML1khOVZWn/F3POdShU
Ef0L4if2J1Pz5B+Dbe4mUAcA9pTUWjdBzDYwweBWV5z7gwNbHeCia+3tzipxNDkAXiESkBQmJL/e
Tw1fQ9+Ns/aRK2U94Tq16FtVuK85TEV2Q5d8pWth7Yo++Sm68maH5YRQFL1ZsivU7fxt8d0End5u
M7u8Kej8QA64NiZ3vVsTUY4lQo8tEbo47ErkomSMTqdD2oCyR1qVoLQ1GgoxGKN5nMY3lrlu4sMK
RPOoAMDHy1gByfMJmrNHVC/w7k3+5pEGUyEyn2jrOjARHd9wUl6cPDvwBJjiH3ssqa+j4tvLw2pZ
H92T/Wjh32uUJQrqmkwvsvtKkN6+6tUtVanL/U308QvkMVox6w/Kd/jvEy3KvWLaqP2+f50AAVj5
0ZI5M8jH4nsFBkHSwZJft07axKTx3pcB7JHKpQnQvKnIN2XcphDPE+z47q1Mm+v4i5hpvu4rZ6/z
RqDsxFftEO0LKNX682IF3zXezFjF1fC88QZNA+9cY9RMmFyZvpB4DsAEKrHe6sxy95TVAaOPYm76
1Oli6WRkjBT7tQ3mI7kDG8fUtB5RqkYwjHT0mxr9vCPbP52F/T2J7UBCsd8Hxq+tMD8+bSgvjo4W
FnTZEM3FwFyan0ljhRq/WwwzYi6d2AKbdYaHwuWTfLBb3ymDdOuYWQfNQmPLCzUNVEdLcE0DKkOR
7ufv/0mmpIBwXSfRsmDq8sl429E4Nq+qtynsU6Bx+nw5jd3FQO3/Wc8fiLogw1lztcT5O4yy0J55
QD17yvZ0pWn8wiKNiV0iFKSsTIibuv4fVfL+gcPAUxL9cqzcZYQrJ4i4FTPc/aLHoawStsrT+NNF
W1Vzi/6+FFtEjVthvNEbW335K36RYcTe8eUt4W2ZHFhUjb/Myl8AL62Wn4MiQ4zGsBEkqG8rWLEN
cmbBUFmTRy95Yd0o0wmoojDKS0gm+Wn4XlAl19K9fniPpd+/YGrFC2uHKSxr+F5bbi2wnNsPRXeq
Miu3lTPUtYWCmLH4HFZ6IQOFyXgDyTAZPb7wtkMY7TYuGvJQFCCWog/AGg3a1yTPT/xyq/XEsHRA
YONTtM8ZsejAfRyfLqMjSC/9Nbfga3JvFmqztb/+HeVJlpBr0uUZFDX2tuJIHHZ4168PtsMOM19r
2sWm9XGaeNoxAfDdsg6tgNxJWsFEu6SrZbrylqW0nKXUP+4ES8HVYUzXNXCAbMBSIHEUQ/5TqeRq
fREAvcYV38trmyppfjR5nUvuQhHklGFMUvIZCsD65tjvZnb8jevQLKT4ED2Szi9S7HdIEJqgjDLZ
LGci/UA7WrvXHSMYGK9GijhsP3x0Yo52EfQOGZ7wU91h+1Skyfk2inkasRRMh5jLkbIiqWKZpgSe
4554YIeh80zMiETstV7z7k0sYeTCe2t8wE+lbGDGXxRYH6Dja85TjGqH9IiFbKuoGKBeZmAHhMGE
VnkNgKpSvkkMft0qlloaAf8ZCmIBl318rbvneVy05636eGUbJ9d+sO1DNA5YV3dYBGAZllbEXozs
tr1QQ+0Ewxhnyx1EhyxGdbLtcTt+oGNvhSp2oWBpKNNhNt3qxD2BfsB+w7XZmNBL7qVDMi6dQ5RU
mPYMcaCYcmm3QK4rLn4TYRpCIx74RFdEyUPF16KJ1l00h69Ke61ynU2DIkoJOHLye/UH5vXbknVk
qqxszxAqOFo1kMUoghoCPMw5hvh31YojaEKQl8KYxbWiSa4V1DqkGRs/LUnye6gIG6qySPKmMZIu
DbtuPd3M5tv0zLraaHlDIVVxNhl8K1ForuEvXhPjJB7gnhiNfA1hD+REsyZQYiY3u5vbcYA0dfjg
y6luy8fxfggfxgi7SuGalaSCI+tSxZEvA29o+PbkvM4rQu56lqgEx9RO393g4tNNbA8c6D3cZsSM
4eN+8tHQXVoqtcBkKJevXONo+8KwuTT9UNOjWfeSpnS1M14wyc7YExmjSXIjY48NB3wHqCXh4SWr
fbURuSA3CHx2X8yu2H5PyWeGbvzysNypZ/nPuhRN03ikbVPxqHAviOrbC8rAuDwkVBbTACuMZ3Fk
leIDnw+YQOLrMm5LP23qm3ZFP4oSAq36uLARp8bLxRsHw6m6MZ+zbQBAKaYSLwpubkoJwUEjzXzq
HTHV1U1VC/kPLyjkaLQsz3Nm8dEZIFvyH9yxKgps/E8e2Z9dU49I7VHhfFOD50lgEEjvb03aiZoh
gMSN8Ffk2/6fLe7EIueOFQPAm6348KqblVlDSQwkzKccb23ryDmVU2hqKboJ9wkPli0BIrCvYSbi
dLMl2W23fgCsyxdXYGW4XqAHWqt4avIFU9zWlEfb2nk5DcTMiX7oP/+5eqiQfiXC1TnzMiUIo7E2
1idTSFhoEsJYKp/SNQLECX1i+bgxnD4EXnpmX0kNmO5OQQx2ck/SouiN59nOxsf8LzcHo2hRzFNQ
Po3iGtk19kYCSh2wBWDPIffPk7D2pyywyQS1lbfcFkecYX1w9gu6b6b+C7gEzp1uXdf63gZXKykC
ZsqYxrb8C2BaPvcW4w4qDFbhp+co7ue2NvSZIbBYEoGCH3EozG/ZT8Wj2Xf4Ief6enIkO2cRTODX
RaZg28SJmPqfKeReJwTWX4GHD8DBLgWaIeb52Od4jD0C5Pgqv44DORuURWP6p7wsyMnLznABzDWb
Egp5/KTZOr567aWDAFPVClXYC3eL1v/et7rxButUa9oIQi0u5YU2cbVN+qvvrsKG+cKYbwoc++x6
sATpgVE7ikx+4CKcfU70yszM8fLyKRkM4Rt+8unPTC9HYKkDP152DJkdih7tisbh+glnN7MxEM9L
uWkQGD8b2l3AQ6KtQnsuLckCSJEQe4aj500BoRY9vgTgmHwmjJgBREHennIFxJTKj85M0nQ+KjmK
lZaZMFnKrrBFVbqpALEv7p7MSQnKQ9DLcVT/RSINHwAZ+U/Egg/BCZzIBi5w5MGDxC+g4/JVsaJE
gOVALVn6ZRhArgmVOaLs0MPZa3PXTYH9xvC1kT6y7cyIlbbetg1Jl9q37gtYCE5Y8Rmmu7qxXqQc
PNMgFLOuwAVzv2msrueOLHmowxAVMkR8KcTgInjljgGZ7YsCh23Sh0ZWeWqRzIWEd/UWao87mTBE
Os5XyHW8ebFugWqevLBFDECvcNZ5u+JriQRopTSvGHavPC+adjvb02x1+mnlyS+70Nr2RBqKXEbv
gi6KWv6eS2kYnrzalhGIYQ4luz8ZyUCfxojJJR3YGtWx+ACy/OfRBlGsFefDIgCqEO6pu4dn56ox
RUM0+PGSiaOZ+3kxrXdqkut33+AOYsniXxGFVeQXF3LxxDK8+E7MyGk0wJDVC9CZ9/y1RTQLhjMS
SclsIm7sw1taaBSwo/HPFVlakgVsytk3h6rehxuRZUSkzEN5BpqroPI1eEJqd5gzKDgqxT8GezRy
urqR0SCUjxpyqgMfJKOKvNokcncJtxd7yrpQ+0wNaQx8CKwlyhsEDMj2yOk76jJhITnZvVRoNtye
3HcKj2nJDrSwlWTV+UBJcmwAmZd4eM5qXoMH69+Pnb/KjAw51Fu1HINmYfagfkSgRuyuaEEF/jMF
LIHr3wui+9Me7Fw/Mfw1+U9snq8prAUCzQAHGHARZijniJ0tw+5SMkfYTDIF5W5tq34VnPQlOn9m
KtM+ZdAtjNAdMirVKfVRFTBDR/XP8UFm3jh6Mv+TB/ob3aG10DLNJjJtyfPvb5SlGi1AVakE6e7G
sjd6jq6rlrpe23pPYZACmsHRS7iRny+xY6bvSZEJXy/o8pzZiKsB6ZitcvaB7HKGhiRSHVXJjDDV
S7DZ2QhMHHDdRbZ+Uc/J0heXeFPSjuZditduQmfxNC4asZvP7/JI+5mnKAD+471jq7kh+dzBhnwn
xCmxMK8ytKRLpCeUnt3pwOOTtmxlpFh3ZhouL6T7qug6RuTHSN7amYFObQKCzBNwZ3+o1AHaCvNv
UqzHYgbk9KsC4T5w4wRozIvRrDk8pOlo9QmaHREvbEq7pc9zMwl0sC4zEht3oAvnHMaNHfwW6yqV
grxcTp/8i+zuXj0FT0ZeumtE3CLlAeInCMUL8zKbKdaI916fN56iouHuJGg4ue3/ahdyLoutBJe0
YO9drc4lbsnE2q11nuU9vzObFIc9QmTX7LYZUjBorxaYvuOyc0phglIxI5+dB2p9r8XtD9Y5XVvs
k/aTzZcS49rERqmkWw//4vX69LmhRwAdTwpeUkFGFCJfecY8iaibOETmSTNTm66jJd++v/WzetO+
wJJQkSKp+iwn7eSMLbo7qTOA7neZUs+wz88d3AN4ydcVEU1MpbCCFPok63p3NTO83SNp47y6UIQh
Z0ENIPk6qnCZlQwengKwS1rD/gDmVX4vipRCBpVpugNxBqrxkyUIoV3de7RcBKaT+mW//K7nu0j0
sTaOL59Z9eNDHFKwokIGk7OAvYccg09eVZN102pVj0SRK3Hl/uKJvC+4h2E8hQzoh0iJEoNk0658
8GAC9NajTOK7iWnHwL4RwKWpgyO0qaJ/U1zaSiHsbqAZQkic/WBhkCXuoqFh0V4LeJcPn5SNG63b
h5EkOiEQWgEjHa7A+rJ0StQ9wwoYY2uelIsoYFAiNmkvDtanW3lVXXUfPEhGiJD1b93UXZqWGeDw
aifzddo/xMKc6QJdj5iQ+AoQhBP2lZ4wriaZylWCqpVYPXXHuFtOMhK8XkkBYhuOUgZi0IOLXzRS
J6XeETkYYz0WhJB/1k1Xwi74QLtAGQhXydOwCdSQejkYk4PLpB0JCgYvPK8/2W//zpiGErdO/rgB
gltLAMgi1F45VLX2M0fPf990dcLusW+8SRYqSVg58lyu9d9+bJedzR/QTbED4SIf06r0wSDkw9qh
kOVSnEr0I53WGeDD5OkUqMqkS1W+j/kyTO3GU16MQVky49xk4/WYagDpba9kLZyZwP0pkEthA7wq
tWBEGYirrdof1PSmeZ3XlLVFyd+PkxluAv8whRQtXVhtRSBV7IU5Rvd4Ii46srBAHy5eJs7kJpJ1
f1/GR76tz9UvVkx2W50rHALwGWkFAMu05/9BK8d037XwXMY0P/8/8jTaAmkEJOVtHhxcM3drIKYo
Lk+ytAICRhMXYGgJXzbA7yqrVr1wh1xBbTbuCWqlZl/67+u1EKWGchkctgeQcPRKeP47mI1weQEF
blRRx1ds+/+XzH4ufTZRMKDI63z0Ewe2LSy82ORjANCooiHocHg00Z6fqWaQz5mOZMCmHOcTl54L
al7d5ksTbPW7iL+VDahEjE0ivSZFoPjuzgZyzw7S9gg/PTfgqxRq6yWcDhHXi2Cn+fwyGwDdNX7h
/Y5U0IH+m15Xb+ZwdrLmbuKGZ7JK0C/l/s/F2p4U5I6bmWzhzsIEMy+Hinj+ET6WzX+XJ3O+s1xH
WnfSUXlPfosQCaueVfFuAAQduPaHjj21l1JVaWYkZ0w0g8HSej6YWoz4JbYqGP+ynOdoqufOFPFr
jROqoZJkGVdo5g2LVwPlw43bksSbm/E1cJBzEOe00CowNiOsDVK5bs4NM3KqNLTZhwWEzoHFcLam
h2P99zrTxIKSsXim+as/D+PPz4mMcjlSBSO+XC8+/y99EC4+RDNoPLJKooLPsSCPUOC+psQ9rEXy
duJef4F7G90zMdSuS4wbeKx5SdTk5dgKhbsE3ReVivKPNMlWr0F5l7/hS+2Jrbcq4E9Ns4QtuimX
A7Ncwdd/TSpdl90jvlfzjmuNDnrn0HqPGoaEYkx84a61YR9mhoIjLB0smCNhsffAIXBfrEl1slPW
n04ZMCUYbMnlM9tqRXxEAgeGHU/jctxOphCxS5OhTG3OmNhKaFS61yL9V/eJswssgLCwOub3l50D
Grti+JZ+jmfLQ1HTQZFsDSvIvjilLNReEuQHVO+47pC72d12OURS1GMH9/zi/2hXs36wP85HqXq2
EQ4xsAqS7RcPgw+d/OxuPxLlmLsIjro3Fn0X+ahWrqNAFSTgNsFH/mxgByHrJB7/jbyeoru9XPx0
/f8eCZDrAhjqwIxGV0h1uYscGwl6A3ZnxNp8ROzP4SJtPwoikLywR1Uy3nYT9PPMHIdd6rvUF5jD
+bnn+DBTuLvQWNJkN0WxCAncDaT0T7R8nzvJ4MziMmEdXGxIecDD3WyU8Cnseq27jJ51hrj239Nw
3ZB8AHIwDpMlm04HNR0w7niluiTNm1ipvjreIqpI1UPT/u6nZPjX9QPIky50THLbWCfY69KsF4ho
ukawJqhH0OGJdtt01ILs24iOZiBG/vLyWqFfYrnO+lzv0eBGRAmrph4Y6bwyetGnq0XwZcg1fyba
SR96kQ4HrvtPh8cqmBGo6SA3xkbK0DRaaywA1TGcK87mTmTG/A/eXPtMCpxhsdOgWyGrkIpdYanH
3B9S4uL9y8cC72M5/beRqCUTDJpYfTxaKKVtAXm6a3gSwxwYKMKerWnp3I8DxoGjInMj6HeFRrQg
P7MEKsRKmLdhjrPvjEOrYetgWXXJnschDzx7WuWz2mSGdsYg3iobZZE1+5VuGleHY92oir6q3d4w
G3uXyZYck1O38n6yUKPDyr8UpslsDooLdM99RjsND+jk2tspvDvXIQvpiOzsaY9JF+I3DvgWepHh
9LMfju90Zl8jW8Hu9Q+6gMS1ap4V9g9WfAwHfarbFKP+kB3eTNkrwxdZX+WR4m0l/vqfr5V7PPvR
jApLikjNK0fnd/cCfoOiWMfk7SwVBol6F7oD8/hqJrcvT0Zwtx6G5V7S/AUZiTT1p/kn/PT9aBrX
whrvrl1RPzcP+FyzP7pbc3wSCu55iM209H+qhjICyn5xqZ2w18/m99ZD6KXfUkge0E6z/rGGSJ/+
IKrJ5WdS4ReTz9/jZGXRkkhKe4MI1CvBPlKrS4VqaBLcTDXX8t78vMFgbwMti6GWTId+iLMhuigy
Ceq8fO7j1mFIEEWIe2HNvaHF3xWmSgyok93sx89ARx1OhSKKtRYc13tZU0pH2MH8ige12coYtuU6
JqgHG4UpSTMrjyU2E4KBBE4YxF5eEkqZvhLuKnHWAL0X7gTF9Uqw5YTWPkWqwp2eIXicOoporceN
+Vmo6fY/YhPFx342Key/inNwH+XSIXLb/JYZ5agwhT/zTodOtJF3DQP5KjwBEkILSPo5nEk60o1f
wbZhOB4HTF84YnY4yg88XKqhjMYx5qHFMMvey1L2so/+rIS2fYzegs3VYmbR23olwq3r5HspG1C7
uIkVkylhQ4bfkImDXUJ977XTpecFSQKO6G6bHjvjrbCHaQYEmn3IdoDS81v1yvZYE1FdPLJCVIH1
gnDE6nHi4TGSZc5TAyS4zCT3aSI4yNBPbLPWMBtKW44g+lbPWEfH1sgA8b/CQFx7trznoO5tJFmp
E9tt+5vyfU03iKNamsT2+3mLE8V9XKoBVdCHVPjOLgEi9iJBIlUPXKw5I5k=
`protect end_protected
