-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Ys5iJ52hEnIk0A9J6pIKDjVKIjejZcZvEma6ZL9lun1naQ0gQGA0vaoIxp30+yw9O7jqKl2gbpEt
UoTtd4AAxhC7xDUsHvM7wgd4MeeWcPa7MwRLCooiSwJnio/0IUfqhdV9ZTBHHbI9tKs4Fq2KqL6c
fomYl5B031E4TGe2xaIf5rEwelHUZCB2npdKlp9O8NrA/nTQx09PmFoKosz9EsvRAiEU2sj0XUcn
BYzofEQcG1YTdWLkItJnfh/fOLHqQc3cvjhLVrzljCA3l9Lbfvykn4uvO8D+MKE3UufRHsSXPQJY
70qS24L5Ch0nd2Mbn9gT1I0xaCsr93sOo4DzJg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4288)
`protect data_block
MobS6L5fj2RMl6feDtEFpcMIWVAGdmNAp3MOHbfCQ3VFfALAKFz511eGiL/FTUnTWDY2mjaeXIGy
8PwMTIxyMopmnuAGq6KvYrxM/8Znn8Q7itB7Td9h3N6/cSXJCo0eI7tgELvtOJN8tSTCmia3ZsO3
CYeLgvQZpQkmJYHGK92XBRKEbukBcFTsKN/xgaQ2VAciUrFB2w3NrS0x0ll2pXlvBMYBDjuCSrPy
MNuJnC2Pd3NgF6IhvOlzI9CS4zP1ekiD1LLihlX1cV/lQT8Z2vi5HpvE22Pqd+ViCK1njs6KoLg9
pImEySVXdIE7GBrdqdrokIJmzEn8wRGCwPKteWFyiJ2yaPuTOvro4YbyKmVnSnXfQiBVJ+/GPJkp
qSjuEnali+rW83e3oM2n7+Ifd9VBFXRqlAV0rNZ9LsauBUUXtDzQafUDQ1QcS1IVdZwFG77J1eeb
myEVuHUluKdqVPx8XeRBns+cARvDRlYyEnS7OPkcIccmuL87BJJxGAnhPAPFvCZN7G519Qtc4Lb4
NpYC1tBoSSUQA8DpduMAXk6VyzdW0zA8D5j9nSQ4OehyPZMvsXDv8PPuXUWBglKSpQ0kqSY5hUHr
vzKMx739PouPHDuaFMfxp8n8eRzodxd4rIfSy30xTlvIsWQ9+Gzyc437WYO4WEBF/1tEifbsrhw7
rh/r3tCGi8wy4Br0Y7vGh2Ns14lHAPYW4Pbfwf8B2v2vetidcH7XimcYYI0/4mT3HMXVqWTKZCFH
MZgid6kCVR5BI3o6il7P4C7LfDM4XYZt2GgxA2wYzdJuvzwweIY1AhQuZ5OkNHrzK4Fst7ocMbbW
gkkp9F9Jubb5IaluVvEZ5pDTYGQRnhPosFTIxW9yCJW9ZJt0S/owEQlSg3SXAk+mQsQRLnx8E+eE
5UuUCCITs1ZhYWClXXNxB0JuIT/WhgDr3z42CbnX3IzMNPZgR8MjNY3uiCxATxLRX+6TyFQ2hDvl
z1kSrJ8e5CIImbkr68pPXbIKlHxFzCe1NjAleefcrpZE4hsNLTyFEGVPjoK37STRkPQx0w5ZTRk+
UKRmp2glp3vODsaCODcy4kWhIPvcHJdLDHcTMZJpYAEm157Ve6Lrm1gWegZ21LBrWHTVnW/U68+2
k3Oww3ypy7CNIz+ZL2Lr0UunlafQCmgKjxLxSOKz4xHC8dS532zbmEnOoE/8FHVUUr0nTodCwzfp
GpyHVxdBxjgvMTBkD3HuO6LCjIxvy+e7EwWDovf++U9+WCKv+MocdA7ND7ZNL/HKCV96kEv/9aF3
GJCcuEWqJbFS8JRSLFhkkjyUMR3KTFxFLAIQpBBxF23ClZnh4SWfp3qeP57DD2WDAuwezIMDlZ8f
rFTCxOaT4CkgpQh+rvhby3lcU7SMmOm29xaJJClzzvPIhCKjOTpWQyCB2bp/Rau6/QE8LcIjhA0i
kNCDJUwwY4X+ooL1jU/vx6dMeKc2abIywjD/JoV3ceNSYmlgoeeLeO+LzCKdN4IuxaCKAG+i+/fd
kxFO+v0n5e8X/48WEvvzASzXJWBu9mWAgMBPvETLJRz6cxuEvooy1t2fdAsdgFQsKDigsfWlacz2
gakWfdi9sdVvEJEuAZmizRU3wr15qBOuPqLFEHmoM5/5F+jqXqctsleyZ07HgpzS4G8gHRVfSuPG
m02Y50UF8flqJigHtdkhb7Re/lT7qkzk9w7xesYovTkYzGYbqlRneFIWQhAqiKehHEpxQJuOmxY4
i38hAB2v8vlxSOa51kecMX7UGvZ0a+8N7q2o8iGzZkE2ARH5qA0GyLnOur6gs4yrqu0NLeN2zJEs
16cHJe9MIl7u0llbIF6219POKoExG8syBVZ2mrJScDad9AjsWE55UXwR+S5eSdoyXT9Yp+05QEZS
QIaHD7hH283YVsYXSJEb6YoTlF4643yDugvFUEK5ZeFVY7ntBU8kTMIVoOPMP9JPxps9DwT1HTWF
MR+bWTEdVitQv0cGYZCTq/4moMMyIQtOfnRwhOoSZUzFtJSo0NzVmZEiZ0BLtFGhgskanTU/ha7v
InlzjcBFGgue7RyBsA4yw4faAdux1ZBBcTFVe3dj2+UfHWaVVX/Xvrv3GfZ16JQSZzOf3psDIf01
pJTF9lROkm3KSSrA2OdkiyXO8s86IRWjLmnTqzdwCKmHY8yZ5+0WB8iriy8YGOxYES4yNIg58/f8
WnXnIUDJCWSlDGC4aNGPoK5t9KGE4oUsAxEn676pE+DnoXKps8hsU5xVUZVBY2+HGMUbwaFiJ0Qm
IwSdKQceNDRcmyIJ3a4Ka8VV24e0z1lHzuMA7l4Q723ixp+JHoGrpp1l49Cdsa0cz+Os8YqMb4M3
VE4ZZyO3RlHLnP/ElQ/3wqPUp2mM5joh3F1NnYFotRPRfZYJKWfM5X8G3bfxq/38XT3sGC3HJiME
D7TfN+FB4edfc9d48WTjDFucfCjnsxYSeuTZjfPTbPvVHmdT7GUXPCHkc8b6YLM0YVbd2mHBJ5GW
avBa/UrozjplBoAnfG27AvX8yx3ypWpcFT9IpEvzeGPrd1mkT/Pcq1yHbeXABi+Sj7ZXkTmZlLDh
vDKVy8lAfbYJeUUhrIrxnYMdDiMl73uRidj4v1Kho5UlmKYTtDKR6zpoDhoAIeVRLsfaEzx+USi4
BTb4Ols6RnQ6vDyraKw2x9f0bJPvQmXzyA/JAWbs/3a5pHaEVmdTREWMQ+uYn9bdvLj00UraOtkQ
mdhBQWERCvQt+3J6gB2LZCFuPY4mKhoDVXK0UwF7fSdlNHEZV6xdjrTeL8rhAp/vNrQDsqy456pN
YnfOreNUoFCBBCZuV50pvsq3ShSGrB/fsupRfaLKabNQ4CEApQpqeb3BXPfT/AHlzdHAUEmfiw+D
qEOxFt5FGEId7uM1TZZCHP73QjurzW9NdDyRi8BcMIQlYDcHAb8+1lui4hB6wIY37GXAdwwrY2fA
oUH1f9am8uWbMj+0ISqGEsMPEMIls6kQBOSVCkxnTMnD8mBKbQ3wNKwa1HscP46J6lnmDhf2bgDF
PFRsRXD8tMn9IACtOoCa9I7GmEuxHCMY6djoJqE0ChD2ha33KTontUSUbNNH+wZubf43dZzFWNTM
cQqyJU2xPMPr2N0NxIaMMu3unx+iK66hlSkLsZFYRs+nS77GQjV0Ui5H4u4Y3CSkndYOa6MYu51G
nkKtpNejgpnNirNOwgrlwbPjbc/yUZMbc0U9UCgItifnQ6nf2fEM+F8e0GGks5aAux9Vu6UR8j3D
lcQ8Gas0qxMgsxmml2b85/D/MchhU2I4hknzr6Sze4PgtPFAFI+RxJwFT4CqSJaHMl51FtzSabSK
/eW2TbFrZwhaIIE0THwhEaH5UC+Cm8X0PZPpR2uzE/J2IJwEWT1BAYVphBpIS2KDhnJjQbkzgy9D
pxN6hyhI7DFoZsN/qnpYhWAf99IXj9h2s8GQ6o65m6J1jzAEPHE9+HJ5SpA9FCm0+aIOOs3mtipi
O7aXagYU0gsuiSq9dLrCS48OZtOfynpp+U4/1EUHsQA2v7EZhXNMwGrFHjOOuDbK2mnMEMvO7IAL
7YDabD9LxUQqHMiIIMQvWIsJTz75gFV47x5hRq87JJ+eqOm9s1EDZSBzS6IaOV51BWHAfCT+MOhJ
EpytDhARQf7H8/pNTHmgkiM4+V8SNKw5IfbD84blS7szbaeNZSS/U6XR/rc222MLy4tSCj88KILl
DuUEfUTmyny1HjZs/E9TQJuUOABGmyxA9sf3P3NUZW1dupTgwTAYbm6ukTsKi8nQOvTsCyargp8s
mrjkgsVg/HC8tpwsXv2rgJ37j2Cj1t3wogvWhVjmI4SV8NSVBXqfEEgQ5nuXe+1wzJHr/uWOwsA5
NtS26qVQE4bN03Y0ZCIBoo4ZqMwUbwFWeQuWGbzpHLZ7VTcwc3X1abyDwJK0FVfjZls1LpRZp501
M0jz3UORLtRrJ+cqYf6VOtvU88PmvpmEHeAG7ZRqxPOxcgDYCBwo9O2iXaJ/nNFHGwA9Hs93kZ1c
Uk4+Jqg/MsWk2y6tJM4j/XA7zgJKWF724qwjMb4vmZg/HEbmu9BdOJe99mjti4JJKTM/NWPVl3/i
xbotxS1WH7AMt8SnAngkLz9CSAxYyQnc0QzTF6+4m1cfzSFuLGKoCZW5Yklj8SFICHw85lnvfK51
PGNVuBqoemnWISQdnEe6XApPT7H4I4JRGtR9g1bINtWQgwKjKBXtfLRDxQ832v8FG/B4VJjpfzD3
q2diAq2numrwI4qHEHxRQwPOicXGGGTOfiG6xFq1TNhoe/4dPGpDchb41FARjHxidB16x//tQn/X
JtU27uQdLGADxFGCTy/6hXQd/21R7FrZcEC61gjHx/S43N9QrwwBjHxlZUI2aObdOgQGH3epeCl7
8tpqsWtR0jOttXCYSgaR60cEDFZSsy3DMjqA7fbtBH/hjFgnFbW28XDHqKkEEeG7BqDZRcy8jNS4
NpWp4bP8paC18q/s/8IaKeSLOnxj/51Q0o+iWHKjONhWRqgDgPqGPzEDbZwi3U3exAKlvn7083yV
RF6vnu3T4SOcK2dAAVwg9iyPuLD2jYxKHSIdHlHnVTQ7q3kucivMry1gK7Hd6V422eDmayG1cnqU
bUmUDgo0d16BBegYi6BepNOFOmFjG0tcXcxWtHL+WSyKGqytX1xRc8nX+ouCYyKEdn2StJXwqG3O
C1Qr9988wCbjpvXr1AWEcsj6NKJYcujDbnq0y/70m9q9R7xlUcYnVkB1FRoS6Nn1CT7Qbkxab4d6
cTMLbLbnFV/vFVQ8B6Qm2qQcgoLJE3AnFyCajXn/IMsajEqKH+lJ/iGTrwM/uv9EDSmMt/SCiWh5
gmPz3bsJucF+VIQOWwZyBWtKGgltUgnGMkute0HSbOl02KB+tDpuIA7R6fyQx/zlIi77Bg9H0V02
hhzcnVnyNEI93AgSWVdcLE4WfY0SzG9dist1UU3IMe3JZzo9KKNZ73NVrV/S48xc2hsT3gupXYCu
RARwanctIcXa/M4xI8r4HH24UZW5mUK/oZIw9dMx2b5IFWT3zwOkbdic3qE/XmG3Er0vFZPhGyGt
2r/IyAFy2kXVP0NUH21/hrxfrbGTuxqNM4WnvOIQ0d/S+JYB1jTt8P/jkZ4Yz8Cc6WtIJj5FetuQ
ja7pPBFrOfBKQanjadO66CAbl+Kb36l2AZ9+B9BNB/jG7dPvixyOC69+16CJNGfrvfE/zjxjQBlJ
gR6RQNpZaWARMN+tTHWJqJJB3C5jHWLjRSVth67TiA0uL9hBdfMRQ3Ecx4r+tUdLDpgxgCRDDHJ8
GZHMrySEmMnOY1YDCeFxOefxiOrrcddTNDDQY38CloMM7rylNe2a4mIii8s85fBMm2s1tGS6ygVb
hFyf1SkZ/s/i/5BH60VbTRwkyHbd1RdJK4R++Ea3FctuBqrT89hSIn17+SItYFnWhfOEkszxBUGt
4LHVMOhQt5ahIYIqzk3m8Mq24vdAeZ1h00Qy81CpXyGlC3YDn2LhxImxJXD8KaFK0niUx5/V/IJO
bK/RUx8cNzpj3DAnxujlAwIIlBkaV0H3GS8bqQ+yzLMDkK/g74c/VVwzE7ldHG2tAT6UWESyCBtY
3LuQOGKAb0ryNf/qNBk9d6vRrbO0X7sLSjep775gXZXSUDBLD6qrFM9eJT7Unvzrnj4edTla0osN
xIXbDL+cF6DgMBpBXA==
`protect end_protected
