-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
t0vW6sZjo8gfnxLd/kQ2BOC8xwWereCd8pZhD8dOoGNGopEWY8ZKnj7ohZC9KtesSiERSojZGTbx
wfODRZBByHQ/JIrPD0suFQJXPMZgkj0WcLUS9xnomhIGZPy4ckz4/m91WpsTGVtJphKMAfunQmDh
5EEc71Xhq6Rvh/SneCoo8qyju7pGL9sEq+39HzeE1bqvytE+ftx4xMI5bHtwB9qI8zF6dWsKhSdg
lU3MGMIOlVqfISIeMPKTyzyrSyrMtK9PFg616150l+/kdSKlk9YGEDM8/vU9LHAeV2B7/L1DgErf
FMrGk45QOsj1hNeWe2K0kaR/S/1KT65XZ8PlfA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24768)
`protect data_block
TBcP8sUs94OZ8L0sQPSPnN4BqnIGYgF1jSgVcL3NvMRJUEtvgZVaRirerfrFJO7ZReZNJ1hPgcue
1bbBzwCxIP++IwoaJm1vEt1xcpNq9WDTbIlM7oL2gV7FgihuITszhJ0zEACFvaLc+MdTlOvqM5Br
/LYD+sn+QNO7hAmm+5q2xo4+dt7Wtw31/Z6bAOCBjyTCsrQ7u5JM4bD1JoeH3Ki32225QZYOsElM
wE8D6I0wCGa3HI3M/mQwPlyUtsFYh6TLWZnqmpHZtNUGmqjZynBNRAPBCE/reFJXqDIe+v3vwN4o
rLvnMwZnTezgOktANAFGPqsuBvmycLo2ok0pIbRmAvPVbdy/AwILhXJDHcMtUor5idRLZ1WHeKuN
6jwAc4zdQ33p2IVT/U+b35w7DXFOrjELu8XXLjyfrbkorm4/58Wyx89ZJvpzFouORd7nf+v4Bxhx
RU5ReB+GLFRiIldhELzLCvrEYRvhCoC/lBImCD8LzorJcxFrB8iWseKk/wN56g9rM5iWyh+ecCVL
AKNrxdloSc3WMs8rmSb8x7nTljxKr1Y95H1Mvnrp2xmXNnO6lYaHmHPquWfPaBcaMDYQc6XqMWy7
w9Y1id1ZosAj16BgKn7bxpyGrB+6PUYgZ2hiV9NiUv0JlcudexuA/+GRl+rvbzMhsB9m9xdLnFYJ
JqpeWihwarLCgvMrWNRJvC7HR4IyOCesk3DHh8PtEHd8Pc3ISy608uQ0eoE1rYlzBqVaPw4LqW4y
v0D6zx8ZSRj77xjxLr/uthki8eqn9Cii3bTxKRSXeQj5knwHuZ82NE4yh/OfxmKeztdr9r7OMp+7
lsQccsJ7nbfQ99q7rP0r2w+HYhQnATxELq9isnXBguqWaOrzrvezF8BQYHwBpj/nTLF/i5poyJkp
9tpbAbprtERiWovVZ46M5q5sYczbA+9Ol5CuxaAwWRhPdj9uWcLAMptvbTSagTp+dxydzDXLof1k
jhbBg9mm07Mdv8EkcB+OYfR6cMi9w9ZJiyc8SaZk4g9xsb9OHAubBEDpfgdxBtBI8CF0D8nWmc3p
WvRebtgfZLQ9IIFLGvlvx4jkPm+LOJSlhUI1IoKNXrFJj28JnBMtw36/7HJy9YHDPJGULYmm8yNQ
XBi39X7puQgNBXNtTQdaQhFqH81eztlUhFbbNxieruNBh7yFuZ9I6woTJFVWSTNADI4DQHvkcAwg
k26jtKkhFaN/NUc/TQlSKo7N1oIm7CE0RLi9m8iaE0BHmmIGdUp/7M4WedPHoULoXbvipWPoRMXq
pzcN+jBh197PgSXYgFFtKL8AlJheiH0czigLwVogKOVHQovnVbxkcconqre3x+Ko4abAzQMDdR+1
wavXk5lUXF9/BwN8Uv3+qHsWSxQKbs8ZFBt+1R/U9qyYleuaN7fg+lmII9GjZ+2bIEqhI5xxHVTE
W22EWLf1YFptn1fiieuHOtg3eOeajkpLXKOw3mWfblMikN1QAYuD2a0QVcJkU11ziDU7xJs0D0Kd
B4kUaiUeESQB3EpNOAh09S+89MQZTl6Ck6YscpM7vnrrE8EhkaxLIsZM6ihfN54aCIBqZRNFyq1W
M4ue6ubLHmv6IKjqC+0yTK8AT5HyjV2CQ8cRz+eQeD965qPCEGiPNeR+4JlgN7U+n89a+2i052Ln
5x1qaoCUitNgz91nAOIo7sJjuvyU37XJqsIXaMex4exB2rufBGcyZFDV055SzXq22vwbOJjWn2pS
5sQKFplzFxSHPnuNNv1DKkgGvgZBo10pigXVscLe9CI8QxKM53mJgdGwiJYG+s6eyoqoRRnA7AN8
B2xPQr8AE7xVihJr/sHiZkGxwWEEvsDcKAg4y43TWksmObsY5dl0mlb9xWhdS/QEGjPudYq+1eUW
2/wK2WvL0In7vRWJ8/KFfkIp7zMNiBKEq2lFjXfkvqwDgC8MS1j4U5x/+XW8wLgfBXMBkv4gYsM3
Z1KbX8OvHfeOvQwIw3MBt9Q4fNMZrJx6aqHqMZW05GxX+hgb85PeREAaiJA0k6dkgLrDfmd+kWRs
kxUenS+rw96OX2X+LWZ27JU7hS4gh61Qi9aaKjx6G4TBmjeBBUmXZFbRCVFnm88PEIFdK4fXdURc
JcIwUoQm3Ere+tPpQKbUu6gXCHJcM+5y6yRTMt/NM5IbU2sc3rvYXbMQnuFbX8smxvkI5GBBT5Qx
e76oxLCqsVl7uXW6yHTEkvlPRXfYySyFJf5WBokL8tpjqZWyLEbw37ARYlXfvVMPHyih8Q06+lSK
Lpu7AHbH5eZhFOBLWhJGi9cObWWQ0jHuIzQob5cTE+iAR996IgISnPRIDGVATrNceL+j+oGl2ZpD
dPBqDPDkTPS2oXp9VujAquBRVVrxRzGn2h8sYXOEIL/kof4ldvs1bBDXWv3LZ1yn+6Sx0CsnjPgu
wJXJzrU2shFCiN5y2ExAAHyceSjsoyxtLZvtx18deFa4sBBEZaogVX0Tca5+e4jc/AH9GACj+uSB
2yiQemMw9PKi2sY9XSWh24oQ++b9BaPSrjtutG+M86FIEZHN7ljKY5+4jLmp1x2n6vNXnM5x1AeT
zxroYU6n1NKExn7PBFXEA5V1pqBB8e+9p5kMdQfHIg/mAQEqbv3HLIy6OS2m5ozfoqvh88o0eat6
tRTr6Nu5Y2HNIaovuRjf9IsaK+4Zv4j9LQMFKcpl4oyWnrYpqVML0FWyVmgqdvhPw/vcekN11g1M
SNHns5iYORoZ9Rj8zluqzXSZRuao0yOjPLExfnFe6qIrfBItG25U6xUCWVeZtuuNKlfha3a+Wskq
Npmmm6W+P0ZOp+H2OnOvON5aaPpvmg2mPXtpOGYcT1KGCuGR/paWXulBn+/pG8e0cf3bNDgSPREq
UKg8DfBbBV/X+fzoE24tJQtVZRTKtXYJnvzDm0KWsE5HwXApn2thyCOVvKe+E/UlTLIIzJ1NTYUk
klp1GmRlGZoRZGg4tUeupJC7JFFnJ2+fK24QUJQZt8DOxb8ShzHZ5lL3jFlyjpe47FUYhLgbEmFa
ktUIQhW+ZOAbCCheVa+JBF6iFnKEOA2OSW3Cep9hSgxURcI9GSLquk3+Fz7EYG8psa28wvAZok0j
ZbfoGRhweUYx2BI3yS1jXSU41lpu73hZd4lTnfJBjF7p/B0UdxQHMsZQXhENfIC2nZmYYkbKFscI
G0iAaUu+nGjB2gwfHL9XWCc6jhFBBeGOa7GeHh1Nb4jCFLrDkNsHowNPjCkopEXo4JW6jk6cBUbN
QpncUiS2SjQNrXL7Wg1PGG4tN9HGqrfDPUlHTtk7PAjj27ugMIwGOP9FF+8kgCfJvZQa/XZltMCO
Vxwrt7XjGCcXeYcgBP0QbAIFr3utXoVPMB9JHgAoUih8HYAdMNeGIOFAYdEDlzpFZ6R2ICog3tj8
ke9svP6npZ95TH+aFxlvYxf5zTxNq+C1ERI6TM6nz6iiNGIxV3aoKN6Y/H+N67SuC0qwnbNTtk23
94/MF9oR/Xx1OMrvFJVmPnNyX4QeqUczq6JcK7fdm4d23raVAZzF6JB7OLxAwRBWxN47p4iENURn
Pu6lzTK4JYSMkADEQyndSdBZEtA99pZ4sTMeKrvf2Vo/T7SGc/ouSi/iFm3qD6L4pQN8Pz9/IaUE
Lq39vCUaz+IK+40alhMTPBdgjUoam15Jz9n51Z1Zt2b/H+KzPemphphK3LYronZvsa3518uxb9+1
RO2lV7hrcqPzMU+vFrq/j91t15nb9Dby1Xf7U7P0QYYwp4vNvtlPpJPCHnh3/0O81CS6nAbhMqRO
E6uqGaDfRG4ln015hPi3LYZ39ouqIkrC678YiroSO66Iqydn93QLcPQIXzhzo+iVHfgsC2GO49qo
ne+F+eIhilDcyvGz9drX6thmIqL+Yr7ygxs3DSSVGAi/SE2t/Q+bBjTGpfM4G0307F8jhwexEAGG
sUtG7lUgxcuxtRhVF1ASAtASUvYxteKIuzaDUmrevOz/st2B9WQZEbTaCy9N8UH+QKQVdTNRwGEY
HljCDvNxW8/aEd24xP3eX9WmNuOv6mehBmSMZ1x19HiX5L7i66RD8/vHaucfq9DF1khyGC/4jEAB
cVxameuSZBmueDW1YObTMe2A0U5FQUqgBrhcmX8sKeeJAKtCaRQQ7wOcNq4iPhIqG3qCT81YrQt+
wkb9ydEWQuEatoUdUeFDEiNIubyktM16zcRzUleHIjHhMRZmUHglNW6lyrnTBCtWlr7j5ScC1rOR
VvOjxmA091/cmFKMxyrwUb4OTHu8HpeC1kpOAcC1ouZI+3Gnl+W8KEePOgP9kDhTWDJXskVus9Mc
2agfM5R9I8qwtNm/OSC9CUkJagUALsZdw4Y3iII8R50XkBl3Ah4lMtsVmYn8xwQnuv89XDX2Gs2c
92sru67TQdU/uj+pnm+nzGjdhc3QX2vVu7ry+P35u/8F1OztMd8CI97RUzmtBuZpLCeqZZU2aNUW
bOZTyCWoSh/OYhhjiZtDDynVNOxhhoJ63DQ/hXpmYay5/Q2dDbSwsRiSYa+d+9hWLngHSgDoOATk
1zwCeM0vjuDhBkRVd4zTRwNBeU3T4ZFMaOIxNQYG2Y/jBn/f36U/cG0NnL95WvrWX5Hi2nORende
K19Uh1pBLsB29UDceg0SJ22NtNLeEXbIRuv6U/KVUJmWIJlwFnMVdiWPjs/8hoi1ov/kICAjFSk/
oJghHz/HjFGNW8RpULgxLWmgOFAS5/8I4UQfRRYo3heDBrgJCWenJvJt6VqJ81C1q79Y35c72C75
+DxTWusSLvpB3jG0aNmB3FPXbgd9Pt9q26TD0wsr4FaQ0nvpdUTbxBbFkQZ8b9d+Kg9ffT4msrUl
3cf7LdPK1D7POoVOmXCc9xtelQxS96BtP34UsTsGWZ5I11319nW7FIMJFtwGeP5L8whGIyORt6A1
VaFnPc+I8liZ4X9baeIx5TJ5Js2eZS4csBnzoh8CVK/rRDFkQrB8cYBgupTLQ7A7WhWb51kFMNr+
ttzCHMtMjZDjtRz/uDOVfLsI9rNmbzHkaZHHprHXlEYQKvnfjjnlQ43zI/DRtuaM3HSaTS+6/Qkx
5zmxk7V0RRr9jsO73FWFi/4kKyI4p1w9nqbLtVPDqDDw1bCvpamooMIFSFkJAASOW4NKLNUMFq5l
dvjrxcAApdcfFgBFQMaWFqAdlOnsw5rsLiuvcsE+OFscxuV4e2PJJSa7cNKHxTJDYekVYmed/ob1
V0lO9OALoto+rV5/Eok3y7ZhT/1QOrlGGtML1NOo9S5IOf6k5RWNY0mcwECi31b8Ke0oN8JQC27n
HU4JV+y6B0U0MSIYvjF0dgUgPW+N+Z6CeW+fgmQrbXLscx7MDKiORl63PqltDz/Kwa59nkS/50Qu
iqTbL+hOSEwVd6HL8cF9V93KoglM4opmsFNVsDgpguqYF8runGZS4Ysf7wG2utGLe2MuOlyBulj9
LZaL/MAJGXu4Ln0JPwbLYj5/TdROaFhRqSRjNkJqdId5DzPuVqd29bnm7GwwpJYYiM+EGmBC92YT
V0KVveMf/5aBA5mj4u8rOkbauxfZP4KvPrqcunr74gOnWj0eh4u36ZEa603f/StOvKQvQQPQs4dy
Gu1tocoX0LPgmkJaPDoHTaiGYYGfaiMhCYU0ynQCaTC8iZ1CBlIozUPX/E/K3aWOM5uU0N1bHAv8
uYQVZBnwuG+bUFhopqXs/XdPZDthfmmXH0UU0GIsvdmabPM+YmWe8sZN+a+rcXmsBcqkCMNrd/Vw
srS21Nzoq+1sb1AKyT8Volha9WH7nEvpQ5/tXJ1LHiZp8piOnZ8DQTnWXO3s7IyuJM3PzsINW6b/
WDjhUa7snxl4LDM26YKW/lcJiqq8MmrICcFavrLByziJzogiu5hh8M3+0hR8j4PZ5wATgNsz52ar
KHk/E+hv24p1/0jASFgTjwOtFPBBfY9Tb2HIRv4eR7l51E+t+JhBHDV6O7r6kfGUTqQEguphEDE8
zsG/JIfJU9skzJb/PqzoM5I98BrhHD5akYCDV06CATVp4nhByO2VezX4m0bowB5AU400CncIFCan
9c/OgqEwzFgHyj3zdlGFK2TkfvdN9LfFDaYHl75yh0jUOyTsaNYCUieFjCQlWeEYrffiT8B/JPMt
KRUaRRaquTeXIT5fWN/QfeknU/LHyAKkg19p7eiy1se7cKK4g4jr9GeKQLpQWBOZxl/e9wc2uHPy
xgkU7n/NZA0tMKyBMQKChFI/FO2q+Zo9PgLUs/RUNmvA0GE19SYN+zCdnGNHJDS1m9+w+DCPv8Kb
DofbO7UZ4AHH0Gv4DjHsu+syrV9el/iZgaY9reF7VykauSOJo7cAsl/kHnrrH6TC7AOKtHqWH9wp
LiKK5AG8E5ZxunGMwqdIEDIt8VW1myIxZ8OXnavGhd8ybT46wxnaj0KY3KTinFs3efepbmM5qjLV
pH7drxoUG8cc5z3X6KSj1z7hTOCxt4ED/t41IouzpwHhpYh95M1f5VlNBUKfOjzvw5RpHko4eq9m
nGEWNuriDGbMcZK8aWgXPP8rovrKvE9f77wgdzDagCDLHredPh6dcjy5fLSn7wcZWLoCwlZjptYj
z8fD0d2H10+OcohO6KfWztcsFlciAZRBlEL1Y08oI8UGN/8ccLQkXRNqhVjK1KEMBFrn3hw0CsWA
0hY5U58oTeJGnFaUbi2ZIiuk/v+1DT4a4aeC4ifv8MG0voU/ekEAJRZjTkZlr1FcriWyzE1SfAb6
h+CU3iVJhlRQAy2iZUz40zxCmj+SMiU0hHTTv6OMZLuFE3qPMr9mBfMtud5phXBWC0MBhmkr6DEa
UpmcRQ4wqZlGpRyQEpdnkQFqI/7K1PZ6iLUz2SZ1dZ4Ht5sRADTMMlSmEOrzFfN8NWRGF1GuP1uU
LUQElLYABXfkd63XWspUBr8EaZS7DsVoBvDl67FLzrfrcRxEG7fuULKSk5tBHhNdD8nGGsRDB0BZ
cezx3EhXHbFwvNtQ+t8qEs4V7st9zQoxzM6lE4ioe//z3lRTG3tar+uAZaw2FQVy9GDXrkziqcf3
KWKEMiKXSiXMKqzZzSbPdHgAg6WdrTDDRAp8LMm6PnGoR5kqCzq+gf/UYJPXMNsj7WAQERNVl6JS
qgHDgeKxJzeiaM/1lVCGI5DN4RJvHLYc2W4i0G6OG/KUkXznvQcCxT4lhVnZHXNQ5Sc5xbygRSDR
S+XcTdw0zNnZ8S7TAM+7TlDbTp0rMr3uQ8QHmuMaOutPHGKZt9Hffk1mrb6BzfU2zV4ZHjcEuShe
5NAV/walhBImekMLRW8M5qEyNx+RWy6oO7HlSyFEOmIcq3kkdjoLm0gxWO8bm0p4HfbRUJfkSps/
gSGOTX7WSlcJVnwfmyXToSBtoMjr84eQM1Q/AWDmJxfssZSh+5tAm+lSo7bevHSqnzLUHOnwABP+
aKDnif9RqLa50FgSKgmvZHoT1r4T4zBUz2wxR5iyz0N+I7fXDvY6o/R3M88pDZQtYEaK15EO3B4N
/ix+SSoYn/bnkGT1rs3UVL6DNuaC7fHApcfsJz0vc41AaiR1TnjDbscmJNb/XnJbxeLIjjRvKudU
6rS+w4Pk5Y5G/TCuDzy8s8DW4yJuK7QrleHgbEZoeRoDH+LDdwS2N7Egv5hOxBzMIQrtHUBb6H7h
8fwZPwqW+7CLN6p4WCZ2AO0ZCBs60SUvORd3EWXq2XJ0U3bTTP6mHRGgmLcrbHrh/a1Gtk9dNf3D
6uT30GrLced1hM5viPVPI3SINVVzzgYNd6RLltxSdGokiEZOL3iYXgqlJKeLohD6k3v7Y4kmjki+
rlIHdRF8tsYgNdA0JkTA4bKAaXWhHbmfwSAiu5UKJWCxNddUTCVjDPejI8JOA6O/L+hwuZE4LgBa
JVTRZAoce4ptOkaxvOFn0Ca4r+MBl5wGTGqJb3BxCkR0b//8CNk7bePJPFJLh4BZzZK9SFQN21TE
N5eJmX2WEbHgjBvh2o9P4ZKmLVVNe2df77OUltCtYV6HbqFytXGmV851eOmuRWLIru9SkUfQu1ue
QVisTl/SgqrjE6L6GqR5jra7l6OflolVI6uos5iLREKVkI43kJtfoEpIdBJtPsqxvrBeIavbNGss
SUP6hXzYDrLANmaGD3KXO0LtdKabiYQcM7XN8slGvq9F63/CTHkVkOuzygjVHE0jPMlOoFF25x0a
ScCgRb9/Z84lAqFG/P7MAr7gLFHaWlyAmYzAzAQ4Xou47l028uOzFyOjlTJuFH7hdVvGKqA8Tkwx
ey203Mcx548MkzAWv3ykzGW57w26b5wUAiRAfI8l7mB4EEyRaMP4KJqcaSqBc59s6AoBYcuAxU6g
zw99jilTiEmC2m4dfppCkZv1TOo5oOqf1amaejydxMSEPcM71fHmXq4EuhX/ijtJTF+gA28earHF
phxU7Ek+ujpvhknddaFUS70sNfddNyVNqhwZSC4kfok3BV3+JWxpfWrL8vgfxyq6mPSMKxAhw5Im
SXhJF93mG9symlbBO2OpHdZ6vLUdF2eVc4bBk5c5ukc4mXiQOnM8n2Nxd70pwYUlCg2qrER5Rnoa
w5bUp84GA8TIAZXukQgrVczRFRVWpScP73M/DOVs8FSRV8oKyZK0c4yhf5pbuiy8bXxwSA5TGIcu
xX39dwK7qrAEwBU5fHZ4mo5IIS8yDaczQKYUoUl8vC3qrejEzx+6K8kGNezX9OOkGyhPSkCcQ/b7
gsvFEfRkXyNTDyj6Kt7Wu+OJRUZE0cQhux0Dc11nATKBgCbeu5J/lRJvmWRvSkW1L/s+YSLfn05j
xvEPJbvRYU4SiQqJPTs8f9t91DZ6rcrqxf1MFnJ8EbGN9UAiJ5vDsCYiMAQqs3pdwLUrnXnJQpIP
AuLc5LQAD1KMTJFu6UxMUfwduwXFR3jqBFQXXwCe9nFqFYSRQtPHE3hi01+PNr0oVnnsmdFjnkw1
epuJ49IHWwyN5fdz3v0mURShxLG+d1IyjFWDnbPcjMeG7tb1+Z3RGujSH9tHJWzhBwmS/lgKyEeH
yMJLllrLCIV6LG1h5HesQSSukypD8bKQFHfx1KjLfN1x4eVXYgTq1GfuQPyUcWgkxMje+/s7Sw4E
Pzl8hNoHwMLEIeLqXYGqMCP+eN21kx44wGanueIpKZRObULrGSjf6WIIBY9WPU8oKBLx7cuC+fK9
zSemFkP406PL4rivrb9g8BM+6pOGSn/m8Z04BUIpZt2ceuCoGNQ9yZD2AEZPlZN5vSic38JeW44U
fascDEDLpKEm9HY77LnMf6k1wYA4Ky4DtMp+lFUe+jEbcTmsGz6UdQfoVUyLVVP0AlapI5QtK4Je
x/V02jPVVVO9r8WK8yLOQD0mz37XUftMiJMAPIp72W+kySoHd73R1gMGOXjQon/npn1X5c44leBh
Vl7GCtE1BlvhYlkKWiSZoH64+0wUb1L3YcIj0oItkv5XGrYKCrPJyMxZSg5DftxueWkP+Jr+q7dH
Jp+PrkYPyfZTZT+LcxsGhx6soEhum+FU74Fwq0MrLW+0bxEa1D80naTxQ6dgXbY7SKc7S5R74RLF
o5UAKllZiD9NIHUFkk0+Ai/Gk0Q+6wE/Km1fVgM9iYfp8vq08SQT2rdPR31Cs7F/n4iEJZPpv/4U
k5PDywQVUDDgZGeK7ATogoWPaIkvmmIt/t64fL9HLTDfAz9EINYuLK49dDBekWzl4uStHU8Ov9k6
feNkYDm+vpDNQcZZymKrx4O6zjJfmxzprMz541jicbBhTDhTr8IcA3Pf1dROcMytguZfqxLW1hzJ
OOIegZ2mwnBKRjOYpIBa3Bog5iTEJXdZ/r2qi0PpUgOGc4YLuzMbOyA3u8uPEQ/zuatJXM864hLj
rhoiiAaDkrUgqL1MrF9y2RD7lcawzpMTWQsFuDPP3LtbXbiI10M7j5qZCSq4UeWGf9nqMYPs2w4Z
SKlFpzYq004J4j9KcJAr3LTNFJ7nFSAzz019cHWAmlnmrcvw2jUYdKl0bCqZVWGWyyTfH9hdndPX
oXa2shgelc7FpM5+jrgfNio5JFFKXz9NzlCJRcusNGAs+hJNr0t2UtVxF4n/06D/PNeV4QSysX8T
W1H9gM/rZjr5WQs1tqermW8/HWkor51y9R0KeWRGY7iJ5VU5IgOVypJ86zGFZljDxUSRXvTqYopU
HT4jy3MMDpTYYNGDPGtiYf5x1IZMd5526KpgHw51ik+UktQ+FEswIt4EWyJsGZOLfkLkDjPJggG3
cIMrvfIiFTZrgDL0Xu9NF+3oMFNhD7JiX4j4365kMg48eVPrm9Z96tnWZqSSGR8IzQTadBbwBpDR
skYcYcY1EpASFBlTYFZdy5CEIE8DzG1GahFQ+JtbFuSrkUhlE2J6jJLOH4rVPOYZcp3mROY3q2Es
PAxN+zlWQweuAblA6N/G71PRr4ECi7uHCvo15LVhXjnn6N7tcP2scbwyFLBnRLRT/WL9c7o/Lvp5
gSIYqGg4gfP1vNfpR6N2daZD+iM5sQkG+74himwALbuN6kILrTvSqjsXrBc83YNJ4a9aezLJISzq
w3v+OiLP4f56D/GsVa5vUT+8Q4gyVc9x+Uaa01x0c+wkF7+uVEkXotIe4MQXxW4B7xY04b8iPWHQ
imYWjGxJfmoPVPPOSq7+rNyFIh3m7RxRQBpumkIpVxhW3Y9jcdI1TaX38BZOiLSRGu8lehN3aiBP
1y0k5XaOnqfe2dIxiaDR99PLDn1k5op4T2bREtnr4lB7oGvVadPUV7ouvrljT6k1jq5Gss2nZFvg
7Hm3fRc9mPCSxv0IgAIQXZp2IfYJpxG+6DFGcUiyYG3yzAC1lnI2yAESgtjxlHkvlxD4gbRy1fIO
r3vONWTDnRHS6HPyrPDihqhyt49H9Y4hXce8xQwXPL09qhHkHz4TN1dcdyfXzfeVHOGa9duE6ScT
2vhp60n2+EZErwBxHpCu6Uoo+BTRLjGd9gzUe0dNc6eTyNaHc30tM9eRa5BcRmp1ooQWcXwmo/lr
iNtHTkGKmjY/31E1raYzjYqtWGH8S9q/G7h0VLBJoa1pSB0dCRH7CbfJbAtfHmnEH+vquNlIrO++
mnhMsoekY+mMYy6diLy3qf9/zAVybC9Io3aZjQDcXAyPzZgztFCUDnIv+JegpFtrh7hcscRFF8H+
ujVwc3BvnXS7EYVZMy2L7i2u3B4N1rSHJEdGlZmQpVl4PgscqcGlWEDiUI5lzOEEXQHAhq/1kDTv
ySY1lBeto7pylQxHO+myyeTMtCZms4bnuAMzvsVNJb5VG8Vj77lKPMu9jJKQ5jKosYMVGapmXuFt
8Xmww3+jQ1yw3PSo8qSJLOYl3rnhx2+S6gJNZ2OMHdIB7paOjsXPRjWNBpe+XbQDcTd37s4j8SXJ
t8ZoMeSWkVkc/bZGqBCLuPYZAZEBj4jtUiJetpUvCf73iISWJD+Xxi3jGanl9c6aihcPh7yxRx5a
j8wQnqmEIf/tGV1P/s20x7wg0R1ajcGoj0ge7C9baXrClA9Qhdg4oz0D+mw4nItp7/bi8igqFHXq
vU1a+3r4WnLbM93ltWQdJhPf0qvjfISurmIjMbk+s5Qjk+CMG95TOe9cGriDMpntN91BLz+k5dPq
VgrrwvV588NrijXLv/idlpyQGtoqBjYctkWb401ZFka7tnMqX+CJMGIxs0pRQc6A8o+XC3M6Ck4p
PehPxakd7zmA11tT0LtIrxAZalOyXJby+jqMOjWS5uLUxDrf1yOIkAPbo9DGiwZR+4cOSA1CQwxS
RzzU4/NP/dwQVT8WWDLispJarjXfvrNxcz9dCTP4OxSVsYsEEqhuyjJHR1NLBo+7dpRolmFfc6YE
piNcYZyyLjWv36Ix1I9nnpy+kO/javM0KLDmBk9tC7DzCyOScqK5BhSLrern1TLIB0TEqnLcoino
JC93HAdMim2wxeA8oK25nb6nCKFjS6yDreLHhLzfLMk5jcJ5zzR6EXcFe1GJulyZJDxqqyK3qwLG
tMZafowW2SSnxbEpeUmlpRC36wwT3+YmfWpUpBYJ66Fn/h6fLDN8Z5DW3fHik9mP11yZkXZn7vlY
tMwi21wkp2+92KX/WRP3ewnpQlp/WhlCU1f2QISM1M4IP2YO/QteoGaAw/baXFDyhDWUAupj6W04
Y2rF/VIpPED4Y6Tpdr5acs+Ar6Jc8VY/2gg+EGmb8sgBJ9yhyfpytQgI6lOaOX10Y1INBhO1z1YT
mdS+I5Im+ZzZhUFuiuq+cnUGEfxd9EWGhLc29zoVe7OM3Yuockl99AqGafHvxauaquXxYa16uKCf
gVQMoQUSTG+UUz6cVD4cobqxsoGOrV7ZxKTSGcaBHyTs90TyDTazt9NE5sGR7izL6YHG6HD/X7p+
KhQoex0zk4nMlXwemFdZ+opSJDQKzWKkKsHCGF+DUFDYopiS8XjbiJRHd0YisSTzbZGTEFlE84q5
f5i3oHSDFy2emPEL2As84Qm4ot7/9IYpkQFCv9asOLuVWnRqdY6CScCRNx9XS9hfTahw4jf0jRjN
NvwwAQTM5e9DKCsQXMptKO02whAk+wPVOuPMbE5Cuwqlv2dDO6RYebZX4UIt5ApmakzXqKOkpyjU
r7yJX6wVXdx1kAsU9IoVRLFgRODaz9pGesR5bZWQeRipNseqwDa+5Nl+0PasCuQ2gI4opD22kcS7
i90tQZR8uc4pqv9DW6QCfwfsuI6XW428ZserwYOT8/wopbMYdco7bWnsEpa17mU99Ots/xHxfVHa
4SbeXl7KHOslAMw4UWKUFxaQGa3yVZSy3UKcZPCV66IgOLB/6/ymgW6UyqNOyYqKYVLiFdcySWwb
Uig5On6mLkINhl24r0sl3vj8Q3xXOnDIU0wG+ArFuU1jK+HO0CmTNx4j8yU9S53+kLlOBCnEuL8C
ZCPMMG22k7qI0OHxGpLjWzkclujb5/ToMopSHRX+LO+AJRbFBCg1ogBeP8Aq3FGuOyXhgXFXdN93
5e82XABa2o5886+yNa3rf3lyy/iJTuDWy/q1+8P5L8VqnMsGXRXw86ovzc8Nu87L866oOj5kC7Xl
nuKrCXCVfDSPGLXbQFtoiAMTFOeIN8rwCaXqB2zAvyY7E/BERdPB8SoGpFUIbppytHlvZzWZwf3j
lpD+4aSJQEbnF/xvTvaTvm0tnTY/yztVuJndmw0ZBZMw08Fe0PKGbHrKN+7JNVZtITNZWshXX6Rx
N96MGLNg10yD1atCxLNA/Qpj5u4pGU2i6NTJyY7rKXqkQ9RICYU5L22cXYEULd0Gm20Oy6+aQVf4
hnLm/J6Ytt/wneQVzu9hhk2QJ9kR1PskYmPRivG0EcfAbybvw/BMWixuo3WvMNZD1I4HYDEa4ytC
vBf75mFNvWz6OphSeEZ23NS4yFsMJxVJLZ07k32C/Z0q3Gdj7JHLySwDjg7T1qGS6U2yRr+LTv6e
UXhqMl31ra2RqkchC2iNZFmxODrV6CgVxav3whgYYMrxp06RitEdZVR4qknod0BMA1kG2D6ZM1bA
ugxp8flEwCpYyL5F/qSp7DB0/zNgubc4ry3IQeMLqqLVPV0P23RLvrao75+SnS33t4Q0rouQUOO/
ikJeN4RI6O/Q/oWY1lhHV1VjhbJ97Bf1d2uUu6EIToI/LHS9cgFDhsUz3gICqWX+HcEXTn6QKsm9
Fb50Lef5/2HYtfcXOS6XAaIyoxdNyrPKLJv7RsgsztrSYg/wuDTdC+MePTrkHwxB0xtI1zCga9JA
szvUypIby2cdBR6w01QgQZVy/BhSR49J52/kEibIsO/TyZ6J6hac0q6g3sdAEpwXMilKWmf0W2Ia
b8UbpHMOsgUVSdqMJN/UzmigfBcyVRWE4Px/gIj69Jcpu+5TLKHM19D3TA18uSAFVGFB1nn5zkR5
BXzhXIdeQiS5+CQeZRSYweAlgwCTg5lfcAboT2yELlmtA17nmEcEwvYX6E2BVrdnK8JYJ1Aw3oOj
8EFW0GOOUnJPEifwhVrIzoLXGOFm/YGtUSco9UMKlQazUi/itLPhcQnMBGSA6zldejdCjHwvq284
ANC77sUy0XOc3mk68UiKGD8ufjZVSVbpNJ0+ZTEJUL7rg2yBr3b76rZqxHN0h6vp50dyV8b8OTnY
tdMxSug29Fhsv2x94NVJVG4eEdElQHV49YzDFnnCmij4xkGIFRcr7hlrGLXSbSvYYY4B7LO7vCXg
v7X6PeXm/FYvLWbv/f3Fhl41Peea7FHJ6qsKtZ4a8zE/Bhiliuor3HcIemC7VzZ4YlcZAbs09WA0
DwRwa6aMcsH4Hit67hUp8S7HVA24fI8nRsdZCU60kREtU2obiHL9mIZVpC8NUGQ/lD6HtADlI6gI
XcBam34br4Qc8vOLjqyoatkVdCkFh4lJvjWku2KYZNJVvEwpDvGXHjl8txyPmi+n56ID7DnTrTVh
weyfnpsFqGT9CMeP2nO5Gz3UZvamA331VzDCd8t4OKUfLOkTYN0Fbf/MRnH4PQP0KKl8OC8f1OWJ
qX4dOwMwfjG6RWOQNAeaZUYQZKMZzItABYm8x4gIjMGvo9HB2hhi8hCOe9EcArHOdbK1pSIQVTBk
gusEBSQx+TihCVzfCicw0TkrEl1i6s2kP/GlXV0EfAyBtdhB5DtsVlnc/aeSwAYs1Rf74RFOCBKL
7HAV5WE+Oavet/uQbfqCHR3yB7SEsTU1uol4bsKiIzNCXbJN7oSylitTGQTvnTTbdjVynVswuKfp
N52nrvaBXorEoVGJClQ6aURQz7j+UO0KQEpdK6A2XgTuv6eOwEky4toNgIuSKy/f04u6wBQI5wbH
ikQ+vdz/PsQtIyrI6M+qnQrzzPqvAuQme4AaLRxZmIDY0HqR0aMA2XoqJpOQcJoyDafBh+knpREo
adfiZHI8QXXvV7Se5hMrmSO/Z4x8X6LBVH+epU3p1PkZJlGPjSj1W3NgRhyAPMk44pWHDo5Yua3F
83XwkKAh6RNXaIHnlbAHH/hGpW0/d7Vp31uoDxLaqfGXZSRMieUELsyAtzaS6Frf2IwBxL+UycPt
MHWJBHlkMEAv0Y8MAxEjSw6OuRSD7GBkDKfDC4igvAI7Asf7roH3khIxTbRpDQUVRoG4/FgbAzh/
QGaTFvt4A05nRpzMBj4qJk1Ai3FMb9FopCTzCexJBQz9fdbdCmfqZodATUBMGtwlvXmrAhmT0A1j
3nWnc0QT97nbttNFAPMJzhF/sdB5FmTwgYQnEm5SCMJX4y56PUq+jVd3QLHulB7KgDcxAoC6tk7L
OVyB/Hg5QgEE3sf9X2tfFirIeXyVHcEiNu2RHSgev6raiOM5prWATqnlPvQwRjc5Evj9Ul8M110u
SnffpbyG55Nfp9oYIxEZFDRXPc1c0HhvpORA74HlOcMXnDg2GnzwKmrV4rFz/fJjzPsOVd2cj6kK
DPbZs5YSUHRYypNLqDWNUyvr1kiQ8FvKM4ECxkWFgrCzYmdSr7VCwQh1TKGvs9ZXHKUVRJiDm3ST
WXD1pPSAfkwf1VNVB02wgM1hgzBd9gqA1aOR39DlcJGCKCzHDIrk6mpBFcv77MGPZdZ4HInbfejB
VRZk7RyZrgzALNjR2eI6UIquIvSZi0eL5A4jyLpCVofEuu/w714nqc/0JYTQjIsT0Vd8I6uYzPFP
EmmldkdSg4+N0leyfVZAfTdxIGeMXbQSdkljvE8oXnHiC5a2tRaBVzE4eHaGVxt0607+BUOO0YE3
AmIV4dHRVRKRALXDtdhyY7hEF0K38IEY0IVQEdfEUqSB1sZPzjD+LqNZZqpUeolZDioQovj1GIN0
2YaWiJQKq9sGWrKuJ9voNe3XbOitLX1pOU6LBqHWY6KWozHAh9+Qr4iGaOQ8+ZMzXBZ1wx0/IZSG
ZM9Lowabyn4FHMK6OqeC8QpU4F3QQh2d2HwXdd3AlvhCaATK3i+qjRN98VOf1Zzbu8v7pgWI7T+z
HLnd+DJ9QDXe3/7uCT9X1UyfDmcflqqIwRi0ZAweA41MfhVtECt/oIXc2zVJPpyqUyHwHePDrjjr
66CyHcKjjJqNP+Fdat8f+Jf50t3Ad5iv6B/upXNCrxqVg9wdTl1DHpcarme2vtpIJETUAUcTwcO/
RytKfTNUM40HXDJREpPD3YOrIVhpTIlDQAhX4/eLIpItODGRDirB26UFrT1jdD67AeTY4hB7NBiq
zI9yYOGoQtIyhINJWor96WjZoBRNPyCIwI+uBjcrPl3+kcMJ1iWqJpZwYD17mQ2+6WM6vXwQxqqC
tkbr1JqPgMh9RJHv7opogJGVjcZiv5wyURR0zY1Rm80X6er8VYVTYDxO3IOqhk0vs8PU/DoRw286
aoNkDC4KGa+zBO5icDiZhaVL+71wxOOxdOnOnW2UNtnuvHUsMvpjmZP0j0MbCZXKhKf9myUDylOm
V3578Hchdtu1TD0JHyhZtklYQN5chK2oiVBllYasRugWpSKkLIyD2slUMSJP1ETIQHvUmTbYl+ec
8jCcUeyEwRaOVVnxajTTgRmgoRMF5ICI/D9CV3BWn7MOM/PqnkhJagm2Dh27d4BU4/FMidCMZTUi
zSDAs5NZN2NqmNbjWmFvzQ2rNQoyQoIm275dXgg+kwaB+kdboEgS+dLdYRJzQRjjCCqfuKi85Oqh
Na+bsmjRMYsf2tWR3kI+prXOK4+Ft7ZpyMLN+j00E0pY3eBVEEIGgcAwTqws06E9FarDMPrm1PqS
qdbCLJcE6A0aE88+QlPSe/m4N9hobvgr0Sf/3a0v/DdhT2pt6iMqRqWOMd4miMFDrHgoiUQqY3bf
FTZoKpzdfM5rPPsH5dOesALtSoQmKmUTyVJnLlR+LX6fAAYu17Lw0c7FtPmANqv/myRFtaxyRrj3
0gJuiPlJIGG3G/jX2BlQfqo42HCk5V8+WIENxD5/c9L2iljKCgs6hza+4dJRXGRQGI+MTuEkOdyL
1w1f2n2keikfWSDa7lrxjihXMM9dNIIEFTBrWhhSuFnURgEHulSW8K70YY7eSbpWEZI/DN/kEf3m
jSu1gvrJAcIpqg4EZx7J/+zeenNBAfUo54RMjSesWXsrxkDTYpLeS/oEsC4orbPTFkdTNKD4EGb/
pCvA2bLJCjtYkoi31U4AZ3J/3YQE068ukeWjWw7CLuXLyRgqsZ4qzabk6iK++n42hP9w7uFENL4v
O8rSu/TzMa7KSFaIj6+q9MIvH/ndRuS6YCltwbynf7Nfbpl3dEhleuoBUhEKcR2wNJAHhJ+u4Zlz
9q+hsFQ0ToUsj5WLg7kdmZDRnBkXbzRxZ+rlYDpL4rhKZRLWXfe8Dhwg1Q2ItRnKF6J9hbLKSD1F
GlK+l2F0Sj5TG0pEHXgohspRyK1xeYbhxn9LUgNGapvcC+cDgBwzR6Sc8zF09KEpUW0g5gTPf3yX
9eXd66CxtfNEWCqwhS4V8FBHfVoHtFLTu34072YaF4lxVgwO7Hl4HKb7Z9MxbkcnRiiVbUZBGknc
azlBhte4Ysr5j3qKy08WRcsgdprIyPmEOQckvGWwOele8bpjFJYP8sA/6peDP9ifuX4tkkaW5yUI
JgQUTMvsX/Ln1+wtRL2G32psw9SLEj+mZpgdMnyrPVhYfmZcr67RMKgri4/q9DLb+cFveuxNQ2KW
tFnNYKZ5zVe7Gw3uAbBtjmsjSva4ufWkvQ79/pLPOM//76F9nhky1826Tc8XKCovpw4LnoJYbOiW
1Z5ICX6XI+Jxw50Ilta/X3GchYOTwwssKN8SpnsxBPW09Cpv3hmNEx2/0sTDjFYnZNYY7SxdkxiZ
wDdq3Ybw2hvwYJbxhesL+KxPSKSTKVPyV4JlRm1eXuGVpvT3l5V7WU6kELlSzIPOXsn0ubwa60eS
YMM44qBsfRdpR9rSzQ2Pt4BPRZRdo0xXyuysc6I25z11PkmtGk1EzYia3osIuJijgteKoHOCOC7W
tS9FCpxdxUkVh9M2lN5P+PxC2BfX5BQ7Qqmq2s1WMAsbKxRJd3ey8QOGCHTS8jRaovfz7gWD3ONr
H0+6CFESFIzlM/fa25MbdQgXn6m2cV10juEYe5e879a+91O+fgZgbgkxECTaKCMzSVFkyqFD/nlj
0RE1Im8lwxW1lD9UKeF7JAHx5/NAue1fRkUussPaXZ9c/uE9kOAZWh6VCvzAGfHLyT7FEAW/jbhS
66DPNkj642Bk0nMLvyny1nYgIux+jhaa8/G5614C7FOfUUcTzXCN4Yn2oS8561JHfEf5DtZWWXXN
Z5+UMFlpH7Ll2oCSHvVetBgIvMo1O3pNo/WKtqBzsBBEsT+GTfmy7t1jy1tQ/RAxPu77eIdrlN7y
/WVZOcc/gIp57+hECvHbSJAjQt3B9Muh3o0w6PG/SsFvC/tbVXkItSWFEB4btzJqCkCO+7EJcZJ1
uh72lqvDAeocdl7x5VihOH5lXWens1lRXIrQX8Y8QlQ/KN7H9oO/EhCRgN/joU6Ihta878K9wfP0
pcjv5c6Swi6qrIOHe4jHlRl02+6mn3a2MPTKWLNfttpyq1ynT6epjwY9JRBwDucy21kFjlI8aYaM
CMu5uY12VKztAVyegBs/qZlP1nkHQXYl6/TitwWG/EkEDVRe1+LPXLAFYwg80AzIcrEbZLfxknb9
AUSda5yCfjyM7OtwJJJqnbIt52KKnMUEF2E28Gqv3afHybZcxd+MKq5XuoqZTHP0hGyHl3TVf0XW
yVzRGwBCyPnP2oSPGljMk5AlPEnNmE68UmxlOs1jqkUd6A2lw5d7V+NY7ciUhlssuvjTtDKyzFLZ
ujBmRKA7UQ/iLg8iSrbwOwcHvScoP1MaiZqYz6uHCslDRTaI68FUslPQWtKZ3P0Y3aQL9BwFUGu7
axBYPxbIBoPL9fzSNNjYVFOD64ddz6zbpSPGvzoHzUaPIgB2s3q3O3bDlMDcKSNEfzMMlGNP5t1z
26y0ELmqWQNPvfcD2BYlmc61W96rSZsXNzg8kUy0W0m0Gl7rfaQLWryEpWzt0Yul6oUTdoed+10y
uI+8AC57H5Rd+egC5wlDH2B9XTYekBSSdyySXNkl4wUII0NPisihi8DxsMtaLs17ch7P928JJADy
ctxzv6rshNs7F5aEappSMAVf5vS4SYlPYqLzsUPacCTfRS+K8zVEIrnyvGs9zPIqPLkY45zHfnyb
qAmacYY+Va6xEXmyDfW+DgDRnd5C1DEGhz9+Ct/YXJd6KGNex0pG8n1WzAldU0mVLZUmrNp0J9OQ
9Ak4tq7xyc2My8+2F0gX6mQxSt9I151U4yLVj7E68+j0h9wauJrISrA84NvVSkgLUPqSGQ6i7Lsu
jywhJjkWTzeeIhrPpZoobP9EiIPf47KhmqFHiV0mp8ULS8HapK85ji/AxLhtB3sVr/zTFCywh7Bt
yitsVFviWe8RQIlIeK81x5+HFg3iSnjKVMiyncgY7M1P4BMZ11e5qzjEdg/1k71w+V/qADxfqrd3
kAxhSfIv0NIwNw8bg4NWPX78ss7CQj14FCliNC2JMmh+sguVrSwPvkkM6PSk2UQpo7K7xqaRhito
jmZbhOrgZcgdVK1gbl0W9yjrBkP6z3upJzEp1bNmNFH1IKwpQAu0GYQY/QMLLU1rMuoH5FwX4C9b
mqVJHi9RWg1n/VrrUiGpBn5YpmCqpbkxwf2gmPgjGMNWTyDf1xE5vdyD0oiDWmJgqkXFnTuGKmnI
J2Fvk9WeCyzn132t6RfX+kN1dXGWpHtaCZ27SJM77HxJ9GZQjOBAc/yqXV4YcNdEw86Qv2rvZ0y5
yWp9IW/eVH68qFyCghJz/p3wLLxQPBR0j7hHd8RlW8W1ndU6TvtSBcjNavE73wIAL85uCXjH6zQT
bZTYUqC5lME4hhZZtXZKbp7upxrNKYDLdg6T2ERX39FdZ+zNHv73uB4nrz94D8TciGdvs0u5Bipf
f+OSQnmlO90jWzhF//+M0QVJcor7G1twyrsNjPoGfkWF48zmtg0TyvsqVnuflVqrLaiG4Vgpvt90
qM5TAVVMP1Kce70eYxte+IrLzJ+SvWEb+yhBHx+3n2hkVppIadroYipf/HwA2Rn0WKP8BeKHmAh8
HZVJ4lYXQMsOtbgqW4oTNjmRMVbrL8SjDI+uQn98lqSqlvEqzDPTCtkxJORt8K1v9a4NjwFeWQhs
VbwdzmLjpkcmq2zPzl/SMKc39/eSfz1qbV/s8DKq9hGrlCdwKqfm+uWuntTwKukeizz9u1NImfUK
KmeTcHRTAbfgg+O2ZuzOIRKhiGLLwJGMDIA87Mlh/RuHrH/ndQ7XQRpmIAXHlJU+/VYx577eaJRq
W4Ivv0QnZD9CEcbZqwrp3gzCKy4lCVVf08gf50/inD+czC3dzthzAJ8Jr+8RQtH5QoWiJMzw0Hb5
/3850jIDNaYix4lm/MEDBxgHHXV01eD5I0flAchl1K+XoXI7mh2q/oAc6z+3aH2OEe1PJKWhhG0Z
++pP6GZ1sXgNkZ3y5N9PdhNu1Fi45QZF84ueljkIOlH4oD/dH1+7c4rMRDEMr+m/719C+v5JHtq9
kha2qak60B6W1XokVAt/T7wLgVBbHNZvfADGI1vSBAgnGOtjLBujtN9+oqMrj6xfagExlwnXM88O
Vxe1NB6hHjH2DtM0cFveqNVkFlySSctpPsfmC9nCqT20ugJ3R1TqD4PtPFzXk5t202Nq8cHcMXxd
3FD5SNccVViE5SNSD/CGHOWBub0CIy9vb0OmBsfzGFCrDbLDl6Q4s2K/jtwFxJAh2ZHtCGL6gFk4
sU+2iDIXdVAmk0uoeV0uXgfEUDYaMTfU4su7GcF1Y9WH/D6ZycE9AiG/Oad8WYPfMwmrOqS9aF7c
ETUngra1lSa7GliB5WJ2MuZ2hZOAyvzMNpDiklisErGYfH/CXGairkQTtgdhvB1h3pZ6H40xZlBX
oqgFW3GAUG4YPntvseoEVVbln/0iOsXri6/MSPLk11o1gHFz6VYMeeP/NQm0k0qfCuASMoTwx4eS
cNNTicmQRdSoXc2wwN9wl5iSxyh3gFn1QEWRcQNIdLiOPqjlMNA2GBBbCnTf+gTvypA9RzXtukon
3VaHI9aH0/mXrdqp3XcZ4CSvIo15PlM3LFl35ARiAZL/FHPGqm8evgjycVQ1z+yYMkRJEIE50y/t
4V56PDufoCZSOf6lqnNLyVy71WtrOt7QinVjuaJyXXPOky0HpmcONK5ePBKEsvruiNjRwHXlfaPM
WPEYbVwim+hKq6WyS4QLi+f6g442m9kdR1hZ9JLJid2ZXkMyqc9a8R/n1GjAf09Oy9gkWVqM+w8T
hULS9Nc86zYZj0iiNCM3l4qo+WIuYbsSj5y4NoMKh1679hVftTiax85OBY+3NTURgzU2na0STRBb
tlw+MS0m6K/1KkGA8F+ax5DZX1FcM8NEYds++Je74zX6busDihgr9cT2sho/0F2dVjKcvTjZPzrk
OdrQD9g9NMkOvtOJtLyQinoqLtjWpK5YmqSL2v2bRmvGxj0oAz/YigY5UzK7K+EVekOwVDvRIxlw
OFRz81NKwqF02xVh2q+7za0fiV/WjcAMRc8qXgz0VKGA2NnL5e0/ZdT8ihqGv8QnqAFLsTQwFNVg
DG/7e64WXse6ZW5TdXajRB+ckrUef9VoF8CpXCw5MNkth0puuyEdavJYoV99JxGJ/lUdG/4+SaN9
OV76Jp2JYJ4ZwadNCHeg+FpVaGxkmwVKPCkiinMcz740Kda+NhHeLnZeHP7P+Ja4drQOr66FbsDH
HRuDEAxHvTPquH61ZkxPxxc7/OgAILepcxh+kBZIfbod/NL9m+fZb7UDStVPpk+U8aaBgumv/MNx
x1ThJoC0dvlLVXQS5Ymsp5V6GlfreH2cdUJn68IY2k+l4zit5BQsoS3qR9rXxAP+6dIpgThTabo+
3h6aqXPqYmlM7D2k7QngjiA5GtA3ROr81h4Xu4a6gKp45hoAVGBbDCjIQKr73OCdz5LWH6GGKMMS
VYxdXkFSr5bZUU0xXH/HEa3fYEkwZSEOq9Lz/t4jyLSFw3PoWfGe5ecDUlHWCswsKydmAAx7sEYM
hfG9RRG/ikn4/l3208gSjNh0M/ciZ4uJWfYOrXlZ8Pl5fnc81rdi/YFfubTJwvMOl1W80EQwT7eG
fJ5wWAOktP59jTaj99IhtvLX5BAA1ju7GaKKq/G7zyrSdSy9nQQtGhOXISnh2Yq/GXnXm2MKR9K9
1vpeiTH+mejgEvsgQvYdaq+4haoFd+7DznsFsEsyKreyh5gtu2p7Z4KLcBZr3rnb6TmvXQ3Ld106
itB+y+RY9cCDETjgx6t5c3rjdOcCH73HjNZiB68GAkuZecaOEDvH+wTZYiCkXB4C45UbCRrqPWOo
nUC1UMio24s/2/19Wt/59QVjUBDLDnpB/J/0miQZxKtiBDsY3AGTwHRPosL/mwNK+oG3xSsR9JId
ZUEOfTHF7VeuWKzQIFzqqjMyEztHno7Yj6AOP20MnQJ98Q/wCZ6aJ9xCf89ARrbYHKTPL1UijRjS
PYOE8BeJGQEH9s/A+WPA653R4botliZoJfv/834dzd5zPi1Nv/q+kgOBDwL4nVgfbzqCWBSLz81r
mxv3mQMrqLIxZ0Hr+OSzRq2p2Xe/W6EqYOHBgAQUvaIl4g+L7kTt5vUwEeTul3Dvz5E5iCZMwX3n
W6hqHtf7UPTxUO6bgcPiXnwBa+wV78XIwzRYN6X4ZkpPAdELXmd+ZOAH+MdycIjbOeOhjEWrAvXG
2zjxwOBtxkKG/whsK+uuy2095qwpJrFbzIsAJxOxKLkKrllHRQKNypRreqnMDFjM1+FXmYtCEIb+
e/RXGoFk/mSV4l4sLqXBEA/g3FCUZicchnIzt0JaCDo04Cr7NssrmKGblz5K6BOzQMePky7vX8kp
HBVq95p9VkxX+gMOFJgdsySzw+jlMrBRLrQHog0/yPUQoloBE8kAdKWzLZaZaOmRZcL/mM34No80
YX8Xq66kA1jVRTygxcshWvxeWcIp++R+OFBIiO9hXKqm0BUrwtN6b0Eprv1rKSheVqOlv1aGQn9w
/3WtaZYH3XMP0RvYY6TIwW4nrLrBjNrQWJdYm451gBM0KWHUkPA3OgoMq71GMv8B+pHEEKJvwqaY
V6W7h/0suXhOT8CdodHxUoyLjDhPAgWC/V5dFL30qoKfNbbl5X1OfIUWTkUj3HDXJ2V7HlB85JQf
lV7oDajWVHf218dqGN8rmSmSv+IRXODwtMy/RnLvdZJhvBU2BfZlu8ME5jJoFBqU0HafRRkqUmWB
/BJKoHa+6j3KLQ7UeCxysU0oCu3pMccJy3z9G0JdgiyP44v5X0lJwiDaiupYhi28yUpoc8mO4dhE
LTcPyhYPepCXqZSSVNDKBlsyXvaWyV1JAVUA/+GHCmEQVH0Uq3ikwUWry8CgTBVv0O3p7ihtlzES
GQigIcd31ZPjUDgqEEB/M7f6x6i2kkrF+6Z1SZcoN3mbikrrR/puCMZF7hYRPvwU+oeJnYes5hHX
g2FUX7JjBzag1km4HeCJyT1ZNNxvWooJ8ElxUfcS0i/K6SKvUaAHAmFtZRUyXW5TkgvoiYK58kr9
wqdD9PqupsZKgXkFWHPLTx8WiVCAyDvJ+jZ939mE0Diw4UmkmfkqfmMJwF3bo3aXz82zbBTSXEJG
P4q7G1C4q6RzR0dFkq/twugNyzClwqgMGJ15D7HbonD9GZ9jNWgYviLbFOcZwfkjSfpZbhJa9YAU
jMsiRyI0j6BiqCm53Pt2XQ4dBpSPEnaPcqxDm21isszWv7p378STY+BTU1T1iZL/7h2G99HeNA8I
JcCN0uP09ezKIKIOmw+zySAdm5TS1h0KE5Sl1nP1Bl6PDNoAkzXcTzQ7ApkZ5hhqCpM4QVowqWWt
PyMn0SM3Ras1DJ8TBKF+or2iBpx4TyDDAOy1nUbM3PWXWJMouFHdmpZWfgJGK62C5tzeBFjomgiH
n4phnjcPnXNIR9X4e9W4OFiYnKxLzbQNrDbOl00rhkfEYiSufJMSu3YAn6HKtkFldGiacYasWuDU
dTLpptwCR7HIq4o0m8AlaaMmG1ZOwM66kH53WEq/Jv+euG8D/jnSnvJZ+J9nJfk1FFPH2XL2Eijo
oEz4FhOcVXZj7hSWfue4GoG02GFWneR9xeaC2lY5QbvQJK6sMGQNC9i9Wop5AKPUkTc2tQ21/tNv
USZtSwChN5HP/46NM/NjOqhfbjBv/EEAqWvaSmSeartBOT2unHJJAi5hxvHp2wjCx2iLj+vaSox5
eIbul3GOvvQKzrEdmAQCOqaiz6vQvFufMy6ueuOvebxpCnMZfiyeXmsOBY6u1karpbJJKfEci5yY
8zfQPfg32SeGQbBWCPPFOY6bQAtz3WILNVI5mgte75MM4Pj9LBj/6bAZe/qkuepjIHTBkYjjpPIK
tlFhjy7qmB6SIlTbGvatmAWm6w5j4eMC4BoOfN4xSSuJWqW2B4vacn8zcbh1R+LIbDSM+vEBOEm1
eRgg37kTo3Zz73tkqufoK+3uQRbACckNV0UlmmyHX3zYz4dH2JbRycPMRm2B5KAE/+RKz3D5XHKW
nhDQ9w8Mg4hwA9Xr9NF4vh+xhfj1BGQgSnkPZzXGh++Xl7DadKuaWXNiz0tBIi8FPT/XUqBe3F0D
9/ma5jXCrGZU5HvjkXgdO+kL4uh0zOWK7pkFLQe4FBE2bwexvlYBhMvBc3+oi0Iee/rhSKGUmNR7
v+X0XLMIfJKv3LVW1LQwR1StldYLsvjY7IqpWaxOHASNkyI9RXsQDoceN9a5DTuueay5SotPkCRO
rnqOIWj6CPLk615rgjzx6zLhFQUZiqqkz6BR2/rLCpyYQki2e011qzY6MEYLXUrFMMRuWmk8otXb
q21LQ2BMg3UbwpAt7JMld1Uz1bvI0br2IlLiG5XBzzjPCEOoVO+dGT0JfIcwazpXu3Ig/7YSnR+P
C0yxGN+Onv7JrHZQs3B8qz9Crs9hvPHqyz5jcxnt3VHlL2BXoS9sg6zm+4pyMHcCQjEb7e5pjXhl
5tZrGFtw4qqikOTM74ziOvoho8vH5b9NTEaasuzOZboUdtRXR3QC1YQkrmXiceiDCEYIybgPIXrz
xLWn1Qqn0fXC4IRgyepibH1vO7TvP45Yogv7yEb+qdu+dnwrY4C1HeDoGGpgtO2+sj7w+efNBupc
t3o2EUeLd4yBXhaASsStQo2bhtVtILrvEeGg9TcpujVDykn2dSkIhw5E14C+pl2/aJ6nQ0LCr6IP
TUwYekSv7StLhHJC0h+2w9SGIA2NbduZXWBZ85idAme6n9Kr6l+oA3xRrg5eI1LQj3GrseYV2UDM
C2gL2CynRldgDNz7gruBHFWVVsi56LUpPYA+TTzmlsL4GhVEJ75xx5RARruEtSfLC/m5HwQRwGcw
AJIgYDgLQvgi2+cv67j5/PE/gkslrJ42XOPs8uWpzPo/00s3q1yOqnhTP1RhAPvDszfBFldY42pX
PkYZ6lNfrGygSfl6L/QsdzAD1rugxMmjzDzfDNpo9sRzEayryGNrjWf6O4fAMnXaAhvFZN/Hemkc
3PE4RxqlFUU+mTwU2/ggX1rqHqWMD1hSEvoQSpUaexasvuybis79ifHwbcIvhpzWv0FtXkrz8v6+
BmUz3m10jIUI2rLlL3+Rf91fmEqUuZe4Pmsk8j3XrhZrM03comOpMY2ATmokUYBJc4jSrZQvP/cA
A+pQ7cq/pt4uPCGddR8bzSPIsNX8q9Kx8An8ibo36ypqNCBusCoPgRvP/y4+c5b9HwVZK6+Luc2e
oilpwO02mlzxWIxYsXw4DZxSUfV3XRGeKRYi9T4w/Y6FK5bRZ0lBpxVdlW3ELf5DhiTKdvhD5y1V
T8MsFPqJI71VktoZwjmBsS3HJZjf+10SQ2ebKcrNu/d5eZxDsju/bGHe0oGVKK7wAphG/U6XjGRc
qC4Ru0iCyu+91S78dr939lAu8o6zI2RxtWXVAAZ1kVGW2Db5ceFw8z+xYicMSH1xu5XzCTwq7SDS
KybwtFpiT01noS1dulPc5GNssWS6bhfq3a0+QDNJBAUzGBkg0XmZkYeWpyAP29oAWgpi431JFXkV
JHAgmzAE125bBFVyEEEGDs7+eNHrSLbpUBzrzGl8QTQmwgggLKI6hxBL7nC/JB22JYPWMgs1EO/A
T6fn2p+/EG1+DPKhVtw+ClEadLkwsNvHH3Sfq2wAScQMntqrKbMtVtH2juu5kW7h6S1egjHazSRI
MdD1oOUsxRsA4L0FLI7NDhCxmnbni+dC8iZPSgjj4pMq4xpZVNyOyGB4MxTcdGPAcbJ93Cvhj7nM
DMdjy23RHOPUhX6PiRY1k65dI2Gcb2UTBSrfbXkHIlTq9qGD3iGY9+OX74WWYejSgAwbELQhCXgb
c5ddZHh50WzhsDNHqsdCoentdCY/Us7x98SdBbGUAhhT3rfmXgB17rPjbzRTw6UiHgDIHn+njWll
YzSeEOvXnFbSDj+0BxAlWH6Tl+eqEqUBAvR52vA7PHfinQ+ArDJA0CshtNfM2zxH9Q4tzMSnNAR7
EFUWs/V37lNTyb89Ub0q1zYvSLpilS6H49OdqJfl+GieAraX2JP3h9tvqHf19NXWJp/m+t6J8yQc
5gXbrWHfH7YH3OTe/bvBxNhgLp7AdzDu8zrSuPoKFKLKcSsM45WDf/vEpwjS1XKbLmOdZ/bttLP4
vIbbehXFgDB8QDVBuA6r2Ti6+8xJrgE98xxp8jCrWhz9JxA+3nDPZLl8eYnJD8TNFvECQZlCk0jF
gL6Wv9GkpHwBAvgfnXqbYkndHaQ/WyZE/pUOpYtCAYYijrcNWWwGVLNkiEDbrWMo6OQtHqqECWaC
6DGYRVrAAut7cI4KAjZyx6ycTXj6m16WlfIBPW0YIlI1/3eHu1/o/VocTNRPO9SGnUEx1kunKPUl
BE2QYCc+wlvptHqD2eaStZxFaUDKeqRBvTKFeZf8BWcR1k9A1ZE5U+NGIgKhLI7Plu/CS6U5xhyt
jL/eaid5jC4i0NYKJg8rLV2z96sRbndp9PzK40r9NZ/4BmLwrPO3weqGdba2DDE/nvJ5FCHUnQ62
cz6tKCeLkmry+mfYBdjHt8C6qI20OA3hrBSsvChq+EChP6ZcJin4RmDP8AjFDQE01wF4fDB5Z7Zz
328yA+C87cLGMT2susaKZn4WnkHUlDI/5/IDdS45tN9M2mf1add0Av2LaimfaoVwvebDEk6yuR1F
EuA+swizB9lts2kry6HIugBiYkdPMbdg4Lh68Yk9c0To9/sd0m+Od7H2utxb1k5pBxMimyrfkJT2
LMIjxTWOqQfEiIZ59Up8Iu1T32iAt0aMHMc8No+YHZ/ZdtfhqNFKBe0QL+aMhN4vN9Wk3b/aUhD3
zish+DyLpuJMtvybYLo8+sqGqWSjOBZBf35TxOUJO7Yk7p5c4Sv1cLLB9t5CVm2ULtDa4AGp1X9/
o9JKD56rkBRnan/GaIMFAyEyKsXdiQF/0LIntWGley/G+f8b216uNquY9cWXR+oTvfJ8k37Tirfs
PcsZi3GQFmMQiqBV7cVgs0YsbJ/CKzNebAbgyhCl6q0AN/iQVKzOh0DTDCGgk8+ozy+4A/JYpgEi
mOOabNfBQrTvNRXLud/pTnR9Tl0PcxDaEJ6jcB61MpJH03HHNW9Ccg1M2hvmbTIkoAkWLJ0aPNIy
n3hqvTEwwJnk9tyZGSQSJKSwLzkYchd8uV0heeGZKzuWixqmuo+ZNeHmYe1EH/bYNHwtHkCgPcDU
JGq0nnDb11DgbUo0hKljpGwSG4VoCpfZVZqOZeF1M9mmmpBy4Vm/TsFRIgBcHx2gOOqYrxp/5Im0
MQ1pDtF3BVK/4vUv0JhkzwXfvhjbP/xl+QIjwB9p92yDu9CyMSIF7KCxmmpQVYdkY3JLjz6rT8UE
0fDCm7Jx3GRWsRZDm2H668ZRZRSXvmUNsGMxmq3XjTWC0SRZqMcPYp/OImhGyX1Cv7BaR8jDBFW/
opgsuoa7f8r6PCQhWBapz09VvXL0BMZFgL7wuEE7nHzOm0UepiRAT1AjRbXD4LbnWQCqShCvqCYz
aozXTG2AYxIMDi8O6QOn5wnoX3XwjKwFH98EUy5/+3uVdtizP8N8TJQJjdKrkNU8pOi3DwubqNSe
HppxQbIIsA2fU3TUDH4fKGEkpNFIYceFlTZl8c35hg9ITfNBKjFo5WUmRWf+ApVAPgl7xbipWh+z
Kk9L/6DNz4sDnxSsufJa9knuHfCv7WuHIBICMgMOvltfFUM7hi7VtFiu32HGTDh45TpZDZEOnJ6T
88azI8D/E8BqEh77AkcUbNqRCKbklAz5uEXKPmonbraSVp1O4k5ZaC0/W+dISwpp+2ufO3B+MJ4i
+7TGyRAdm2skhLVNz2L7GMJop2EtaYxW958SuizKTo0Zqc/o1MUlJecGsoHkfbDdpROH0mBAXmtN
/ba2o4G3iU2XiEWtFUksfQ8Te8owPyG52MpzNPhSsjqO7hUPohbdIgjuwZc5AXxMaKDdMe2st6si
alIexu2TWrCis+am4vQ0KL7KzB+YBFVMtvKVa9JT7OtCvLoYRHbzKWiCaSFU9xHkOhhp1biI9EiV
jmOeJeSuDHWtfJU3LvKq/+ZbTRvrvpZULIdNq57BBDldK1r9/8P2y0o/eAAPnkzEpCsFrZhMMFwP
Lm5CAgDhX1oGoK49Vx/j9JjcDWGrhXS8qySd7XcVwBnKFCUbSLHO5oY+Lu2ywno5jJY53YbiEjVi
E94W3dbnwYp0EJSFt8b5Fta5Bb1bN70P6nq0wldjWyiprntbf0unzPIAd1JfkW1tFW5cewKCEMUo
8WvzN07wHgpCE+At3SywWU6n14DkrerEc+IfJlE/3yeToc/d8rPzlaXR8svVealf2Sw+SNVlRddZ
bBgpzcr9Gpoydnajf2X2gMxgJLVnYNP/GLhupRi44bMHA+47iXqiiIavFfao4g1c0GHMSESrRER+
vcViIxmzNdZpouvwxNw76PCanQrIGKdZa6uPJv1Q6+WOc7bB9Aj3DzwLgVEGHRj9OG4DgVU4duSe
AwsM6AdliadPbIhXznGxijpludkT5hysedItZisJ5Z12dbTQa7CZA42qzfLCu4bB6Xewtn2/PA2P
wwMhcJ9LYHl+HtCxh3GacXHmvhHSExBKA2e56HlAUW8uJBMxcFRNH2f9Q15MeOOhraZvWrLHVxZ1
COyRzDiMMSZjkH55DKA4+IhLffE0A4I8gvrHet6srAUrMP9DyOzkzEOIe0aQCx+4WfFXrNoy+koP
0KNfYdWaVJ7otsIrQc3XpEX6myscC1J1PPszTmEg1jmRd9jcP26iRkbO5GP2qKCPBj0ZKe8Cthq1
AWnS3To611sVBCBUJAOU2tlkE1tmp97cJd9GPQuP4dr1bP0wqHI3zEVlFiUZnCaISaKoLfrtAwwx
wKFTOnZqqhDoyCTMOhUOSMB9c8Ng//ER9hNUSd2lxFoxLUZxFRqQr8xP9gu4U5yeMjCbrmwyGcaj
SvGFADXTIfDlflcGebgX106HNc/biBl+NmIJFZBEUFlQ2jHoidwVDL/b0kboySwD6931rgdzuDUY
JTzw+Si+V9zoIZgGeNmpHrnmTIxp8OJISBuRzIZ5IJj3TK2YphsMGlxf+mOQ3+/82zjNI1cBG4Yg
NlLBhGejdpHRzchUK3jxMtVP3UOLcgVzjqvy5C92bhN8B2/rndpCtMeFoaYFTEiN2EJhjfqEKV1k
F82l62gBQV4WCWHkEOekGukaEQixBnFoPOi89aSqklqx/Tqv/NyO2xACmSek0EGMfhPQ41VxtMfd
DpbEirb9YAfVOvpUPUziT9QLuc1jBgzYi65j6cmn8KFF2BVGMSaL24U6wehUCcWf5mIjMUJyvEmO
3ld7nV+ht++pq9IWJZZn5KFb3PSUT5VcppcMOWMV3m1PAzWqrOjwTZe/RH7vbsA88VlcNXHH5CHW
pDS4dKFugqhjZQKubRpuHqxv+mCYHwhhExF7+zFu95jSo6QbTd7QgJilfyukKFtb24sE0yXi8/My
R/VKgCQhpJpNPneaVFvTbz0m8lmpttEdleSdR1Wd43z6eRjk/CSNVM0DKOoRQ3lc+ZVm4M6HRM10
JaWMK+zmkCWs1uI/2kYjNWHm/VMvgtICCpZt6Si5SAWRsRjhE90TGjj9i6a+yBeFlN0N4S569bqb
XpbzvtzgOF3wpsi05BYVeIRL1V+2nVXoMprzFV2yIVyNdkyDNFyM55+5/fP2fseJgm9TcRTC9uAQ
/zccjXGiQB4mgJu8MIiNYgE+9hN6sra0UKGRL+z9s2uA2gJab1TW15esFgeTzy1TKPUO3Ns9zuCu
3wqRcXmSmItmc5MPYsJwnxFNs8FWIxKQiTgSc0Yore2U6Dp+70Etk4/ozLF4Ym/PzTajdBdKpR1c
7neeFn9g97sYLTsM6+Qo9PPWnT85LPUraQ9Eka9ALYHpUwoxT2SeeuoQuGD3SH7T4UY0oxpdKhEJ
sfNOo3IDWgxtNPfdGNyXwesjGBK06m2SAtnT8gz8Abgb7Q1VAlJ73SHt6eZmqycj2P3bhNaiuPY9
miqJpAQe2SnJ3NEBeaSfN2ZdH28kpWQrBuPUaPnwFUF8eCYFPCdClh8TbnnVx268lg1ars3t9+Wj
e/gVJW1wC76iH5naP4y/zmUvafX13uKNQ+sGNGdNsp2BhvaqNzdch5QfL9ggB8Os9fgC7hLzuwfw
S+22LeJemPSN0mQHx6GTfMewOfoLfoHD0xvkeOOjqs3sE3Ke5n4G0CFgsqBFVfUMcShOGa2HyURI
Tvv3rLayixEpr83hbCm4D3rY9G/JCGmrlYQDJGZV9jcUXjdwvICwJ2rCqylzKXQxIfgfmsNu5Qtr
HX6QJRATP6WNm8GwUZhaXSagi+nm3Ytwt7cV+elGW+rCY3rTTa5MQ5JugA2stMqWCh//bSvDWWa0
Df92jlBAnWX7DxIBYcATspwOrxM6zcMPaD4pyghw1eYASCT72G4JAF45+vyBTV/oY9Z0c90Z2rcu
69jJFRpUhwn7xm7ZyYzZ9vUwkK7xsekwvUJkrawwNMjpPk+aA5Z0FEQ4FbASTihkkotxHLK5m0fr
2Buovrt1Vy0Mav+YCxrwIEgurEpMpRWzdJRkpDEkft0JjYh9B355xKewaldwBDeGkg5O3KHntn1T
FvR+PMwnnXgHKHNCriJ0gRSLBo3j8yD5gfYwgqQliKILrnWcM8rZyudQVd/uauDM3bY6W7uHP3jP
4LPlTW1UfadRpRDyjqvbh6Ic9X+JJqcCfJD7+Gl7UoNNLXY+4TKwM2eZ+DeDhcIYl//w9FLIp/Yi
h7Qauk8mA775Wa7o/U6dhbFGbNK2xLFBo0a073GMmsg5Hw1s83nCfKKUOy3mbQ9q6F/HTUdBjKoS
UiMJhP5xktzRg1DcZ/l40JrIdUplqq99GxpOn+/11ojYuUhGRean0Emv7ayQmYWOfIbJjeRFJ6z0
elW0vPUUdIhSaX8qXsMI/00L5SdRcSkvbaCUXX9ZbR+8F1vOHrNgMmJr8JzWBqyN5NVo2pOXIcIs
PYDjjKHo4OKOjtCn0TqzGm9c/k5jRfPgTMK9+vCrHHN4Se4cP9/PuJTcCgLBkAYmrWSvu1/oiptd
gurIbcCh9qVeSE5OtfFL8SeVcZkhSzdYQM3XrftfrBC1V1FLJJu+s5aW26eeo/Y0XvRrGZIJIO8n
I9qbKdKSHkqiRob7Ut36pTLgSRTh7Wu/PGd+7p8HkN9qdkh2xsPapED9cR+ozIGtofdgUk7EQfKX
seL9T+RGEXnNMt31QetAgQJuHX/gM/rB8sh1/m8O6Rs0UWn/sEm73t+Qq3iA46iOsDJdE9+qQfW/
QeFGOoiiutFbWMfeAjebHIK45wHQ5aTsRy/SLs7RLjnUd6DDXrQ8l7BK9D5xbT/8mKF3YxCbsBH/
gYwEkBN6dMklqn9HCpFlJhM+zTbvbmvJMWJGNKf2jkpNnIysULWysl8LIlmB2SexcEB5RGvTeO0E
wUOkYj4ZaYzFMnbsgn2h2XDMcg4i0huVVRhT3wdUNEQK/5+ScExIGovnIFkHho9Wz+WDoXvNG8P8
N82pIXiKhiNJbuymBxU+u/IgrzlreNFvKJbXx4gNvn9OhiAtzCvY6FOlpvdmj7g/Z+QSvju2opQN
gsKSKzkhDqbQ0X9Rjl/ISs0VkhT2GNvvpqv3eBVX+PlbflM28KeiOYu6Gn9zvZXf0JQSozMNO53Q
J7PxZ2ZF0Ur0OrRc2b5kxFPjDo1E2HOLBB77tMFsfo/7T9NX+n+88KvWzkNIraylBH2tAGitsjvA
2Qfi/AF89y9OLkT3qgltPH5kqi5Aary6Usvtqmk7L80xISuaS0wCd2cHd5Nd+30pjV8PNPW83ylQ
69M5KjWKPd09eozlJt7AWclITxVQ3SyGyfGM4wv2XYeVkCJocJnXhvmviLXkYGNB4AqZDZy9tb4N
LFp9Yto6OU5/3+wA7unL9swfpljweZjvuks7kpu7ADCJNqNhENwOiy9I+wQn6fHgGDtpFx5iMO+a
f5oZdzW+c8CWmofk0eTF4BJnWWvK0mfh77E6XRymOcrAZF7dlEpm/8iJmNxxHejEEGb0NDkzvGQc
dGWoedCEquVF4mSt21eBnhUferOdfhB3ykP+79abbv/n3H5EHSiwB++pOVcBJAfvXDdSWWrqrWXT
jrJRpAtpo0AApRB0/3RwqV/UUbxxMDMGMiVkeadaaWcbZrO+NNsp8tWfBuI/o5haLfLWtbl+GETV
Stit95g4O07cgQmi2BDaHNXJimblin5j1Ly4+W7qUOBAL2CsqP1ZQqkAGx0t6KhlgiGlXm5fTmec
bGYgrcD6oibFmNe5HdLdGFo2FY1vfMKQp9veSE9WJy9euUyegrPsGJkBU0yqFZhtzf9e3zR/SDHI
5E8fsPsGR9m0s7XSdlKrTH5kkDdCVPxbV5d+2aX7oW8PZ0T1Zct9OXlWosSDkiceBkJIzcK0XWaa
+6lUkjmcWaZfNgpj3xv/Cr7aZjAJ7yuBBaviy3h1
`protect end_protected
