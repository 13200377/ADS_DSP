-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
z+Q8pspE7m1DU8UxwFHGcuBiJIuGL+Xf0oJlMvgwPmPfcva30MiCDyUW4onhO4aBdqGwWGYcxJps
5AIKkwNvLZf3XvRBTqx4dxANLfK7QZTNlbIswfGaXuOm9BSYe8Fi2XMOs39KaJz4snansMtO3rXH
dJmP4KeJL0YjMKChmF05Y0Z2OlrFzmSEhiXHHJ9np9uNyoTm4vCnQi03uDYsgbubSz53UV31JqMy
1XTq0KM94wIoGcgZ7Vm6H1Hp1gV/vTcC3BRqoHyP77QOgbM+5Tbct+6yebGbjGCXWjM6vS9PbEJh
TaGdVgLCvWQXgetkjE3Wy6egV3qHeko/KyF8ew==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3024)
`protect data_block
LwtDiEDNCG6m4SBq3SeRwRS91NPru6B6GK9IvtZ4Ew6WueL2bjPy8iRgJNClalk633wT7ZFImH/X
K8kT3S64IOsHItym/3X5CHprXTBihqDl+UtSyuWnVOHiKcGwpnWYgSvKw+6xCYiYF7yATInH2GnP
aGSeQC82McR+NzAm+hGdo3W0Z8M5mmwPwhCCvsF7L4JeRm1edJnIBomRYYfEww/ZtmnZL9XPUldZ
gB4xOwRgWEUC6t6FjCph+zG0SSdbgJDEbUUPPvVeJd0qdYAS1Wif6G2xBdnah8akxd9ce36sGvhf
uqXbQMUPJ7KwrQdujaJoTM6vA0EaDKA7WGT/oZ1tYnHRApR9Cmx8EIC9WlS6NwWwl5+QBKwdUZ8a
nDDTdqEfKcPyePMDtR2G9J4VZDi2i6Yb/0GXyQ8EM191yPw51IitwL03EwZdCTYejS7kxvGZCESK
vmCLPbmD1vLyHXXZj/d5An/QgFnYcADiDsAkHYDSqZ5dLXkTS9+YYRtc34zxhOz4/LGFSTjPv6TA
KXkq3VOa64Qp3Dvd36KFcVN8WSad+YV1kWCXZX2skWk8XhJb6kI3G0qPJuh3tjox4wwHkJAwv43U
Eva40CH4hmHFYkZNL0m58X3yleOlOFwpQX02VhgWZM773e52/VohbYnujdr5TVYLTHYD73PWWNYp
UX67BAwJDwLxZa+c+6EwPjlUpRWZFig8qjf59WWKMQQ6zcHsV+QbMZlANM4+JYWeomrVvwHMPO5z
jUHnkxBZOC9nQ0v8ywEEeSyt6GthfkjMPFKFBo88q0uWhYOChwtmNkEuGev6Ue26G8/xre+TAyMa
FyNrt9cG8CmTjM58hciUsfGc7f2ND0AuJXUflmwUkdO5t+Cqt4DImZDf4md58wJCJY06YghNXdN5
jaEFLSrCum1SKeUR+iDEWfyPHNSnOOHIXFG0yDunEWEPeLEGzzNsgVweYaJcQhTqTszOpELEF/oC
ptvz1HQciBTO6IKUGKg7lWDw3Mbl/3x5s9Qzo9qIu0FV4xOk3KI0u2tarhfjS2bF8ppMxcih7S8o
TEsHDxXpbrOnIZ3lon+h4bZ4RCLhGhBkTGq9ypLAxdc0vOTB6dGmvkczsGB6Ay6dS9Sf/SyI+6Um
k83jqhv+W6dtsOnM0sGVffwmgA9c2caJ7YE2s5A3LxeGSvPAgY5FGjpo6osQku0w5qGkfr0VQ/Js
c8y4INdYIE2Rer/8Ufxu7Kh6k222JVvn03tCnwEf/oGhYReC4YeaY75M2ie6fQMh48L9Zj90ZB3O
9mrl083s8dFDumX+8ASmvHJWtV8tUKXo9jGkvp3DViybUnbrnKw9c7BBv06lcQWQDf1LytSDXtob
tSfJ6ar/wbD99nNnlfZqUHir+qnoclL+WOQ7gw+tC85+31zeCdplg+BBbgSKGqjv0GXLQEys2O4F
msEnNHPzYtgK2SUBj+Fsa0o4ObQIuKoj/xKGIOJX+tfj/SIfLFxcWSe+3VyMWHachd1KCEGMwPR2
BJ2F8wAHHEfsqtE81wu3q840245U+wLb7CLxBIMBrUEDsQh6Muk4SM9aArFIMq2a/fayLgA31wTs
/CadLT2NHqFMgR06Euho3oebh8e6j94KvPSErV+fH9wFI7MpUC0y/Jn2jhTV8ZCwUe4HgYlaKPD7
vyJJumD/MBJCnXTuTy6aHrvlLAVK4hCs6oUjFkJvoFdz/z0L4cU9O8vCCLSUafBTz7lXcYP3esVD
9znrRWHIFu6kieAfjt92C1dKHtPZlp7L8jzPONNnEOvEWcyNj3QKFnizufLfdS8Bh0n5otpwK3c5
1PowvqggFGXQ8RP7TlCgtaAMyLmg8NAWYN1Qu00DySutp9G1bscVmRQ8ef4E4Qu3op2VMEQWp64q
IJBfGzP1hOWJyHYeVIfqmG512TROWdCFqBImn1YyAfSCozaa/gt4DKsNR53I9UBJlDpDQz0gTwAa
QRHpWjjPIEEt/ai3Bl5tpJsLbfEHB+AWySdBdyhqNzXg1957/Pzgz4HcVEPDjPVwi0SXkTXV0SaG
pwbSnnxhnT8un6htUGvhTZkzVFPfkgts8L65tjrOv4vDnZcMhZw0lcdvVq0UXqRHBDId32Q3grCY
DKxLxu8NyJVVDmBLORhF9xjLkPb1Alxb1U77zlGyhZCKi8D+2SIetgDT1ET+pxpUnrDpGi1KX5/o
sMNm5J3OiNEgIECSrnGIJRXqHCrmNwj2MyWOVcKczEdmXQZyjbspNMYXTzROeG1IINgyIDEfeNKe
Jsp5xX/32QVmuR0ovScJ9paYw4ka1zzNz3T9UX3f1zfar6hvCGDrs2/HJhTF9+2X1mp9b9h234PD
fw2RzSZmsg5biHGkzQ/ED2aMF60ise7juBQCr4elVx/2Htd9X9GTQ4t2Np/VMEDIwrWi0RGXBNUc
9y1irCANnE86kAqk1xx3JdCyqJbngXUKJEbImwAGLTRMT3sTcPg9G9Bn03ZjfdkXrbVE0uBCPe3u
odt/La/Nv4ouucWU05tplBjgRbc5GxJ8Ir1acYbpbKIZ/xdV8v0SVo11f2SrYMtBvtoUf1EKXTcD
BGGFtJNjL/jy653gtnqrsY7WQP/V30iIL63qauWkDBBNCaqjyRrHmKlrktjXNC8yQaCvF8nD7IXO
1f+EHElPxkyYvTuzVN+4x+h5uyVieifi7RPahP4xaHoxAOfjim21jIDEK22UGVYNWr6OCu0Myaz7
tdmsUI6IOVoA1psyICZTIEhUj3L/wRXd24rNhTXBNs7qhJyBcEStZFYlWEU1Aj/GkpYontkBDImp
RL+FUD0tRBj5yF5BtxWt0MOaqv+XPvcaVdWgsPXRW1EHQfCAlh6yJnFPJqpebEaGGAghIN6bMv5W
j13Pm71fxkjyRMS/IZk8E+EvNbzDy7lcPlcWLHYlygiAhxtq4+suKcSfC5QK194L5OnF5T1LbRu6
SNXyfmXByi+6m91Ir9CZERSnlmnaxy0owt5dM9Rok7mKY4VLX/nBZyXmnFNoNS2v9Vu8OtkEz9/6
498I176U6EIep38OJFPY6P5zh0e+5yEKLkn2PWQVFzUgTQiFc/zylNfsSS1qwIbPJy1OmnRsMQ0U
LUoYjRB+t1Ct8LHhaJTM4GFwXgz4zEwXj13DoO4Bo12HMcA6dV+Ql/CfrygcJt+IhffFCaSuwkkh
iFcGoWf3o2SfjAignCW29z4XiEGENU2yVnfimB3sZs4zgL1cyLIN4Hty9oFLPfAmc0/eFv7/GnkV
YOy0K9OQtYfNo4bR1HqmHAvDBBjbGdzzvd95YOEHBEWA5EIo6eJpmAxW6fuTprJ1hXZcNMMUvKYv
9XZ2b6mB/FboFoOjbu61LMqcSH5GmYU80vp70pz3hLSxI5QVEkAjMT7k7r+Ig8GEtyTQE8oVDLZn
kRmkMJ16M8sqnlcBGudF0alwNiBYSepWvzkLEf5B9fTDBouVoF8WGVuUMiTl2reVZzC1PPBN5SWR
O0E/5YrMKRoUVc/aDQDj3u+wx0ytXCTvfjyRM1ONaZF9+xfTIhS61V3IeLWeeVoDN9ML0wHbYJMd
RBMHAcoau1MUFaZ7ctVgJUpsz7tXYFw0YLsMgoxNyVxofbPlbe3SdT/hPKm0Qu+Yq5hqwClv33TM
MqecW2JxOLdiHDB2mFJfAVPhsO/ereYXxLK/TrWR9mNlt6s3NRpavAVvCoAMF2KcB643F3iyL5kB
K25jr7xAam3vQ8F+qyk3et+27XEAaUdZew4VLa/HdaQhrbLt/4dJWaiFwFxT9+l+YdWN1QbnELyZ
UMzqcXRX0baK9FdEt1n0grTI1lJ6FUaYOk8f1R/nxLfncMOQWmsOFVT/Ip7NbMrrM5GRVqqYGMJN
nskny9RPuieOgiRYwtiHmB49nXZOREMEksKE3B+gyLwbb3mjxU2JHtmpSGMLbw+Sgcclz1l+DAcE
Y6wpGXWIODS+W4DRCwzuwyzJhDq2pY7F6o5yqhrcMdgRKQ/WbxpUuFnF87HFlQC0TADN3jd480FO
i5N3
`protect end_protected
