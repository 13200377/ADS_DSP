-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
MbpDTQBQORYO6SU0QhkyIfASCejiGjxOWWBYIQ2ZtbukEb5YxlpNaQ2Av/jf/R77q2bSEz/hfeu7
E3ogjpE4GiE+nvCex9mU+yvt3logHOSaDZaVZc2YaClXRPaSz6LNxksz7j6htYa+s+TRgdDve8OS
bMiWn4XWLM+7pOd1Mzfl4o4eZhGzOw4gt4qZRRQVKRDtN9Z8Noun6OJBwIBzjJkMgZRQkZQzkHrI
RrkD3SDTPbrH1Il+Q0nDu3mpT0rnelHoCrCC3GKOFa2eKtcZLfv9JbY4nlEhO9bOdg6Kl1gCI/Rc
j5p7yU2Do6Mdc5BMHacbBkjfYr129pS86HGzJg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8208)
`protect data_block
4RwKqhKgYY1ESNneAluiVJkr/JrHrxyAq27TvJOiWhzEbpr4Ul1j3FWzARhafNl3d9HBzfAIO+wY
G9OXm9+GcBwCyWRPAQc/BhK++ZYVRejybvIk8V5cSfsVLOI4e4jlkLaKTOMus9b6+E9dFNtlmRER
XThQkuAXUbNvDgNTQE6nGRuE7KfhhrKmdzdWCId1d7UztUU1dmMfGwn7CzEoXqoIJyZpC23HIcA/
VeShVgPUQ+KfDVChkhCm1n82oBO7dnGRMxjFf/sIpFh5bhry/vVrdyHTQYfso+l+kKROzDizPoWZ
mzjDuH2jMIQOfgp86gdiG1uovSCAWrkVXNSSu/P6ipFVGQwWtojlcJjO7bbAIPl3wANYO+AYQtu7
sSvxUbaU7gn+rmlO6pW2tid2XKaBVrtfVLHY30v8D+X4HanCEqA+UHhfq46ALd/M76Fb8COaNomt
i0hwyL8T7dikC96v27x/2PK6OAZKQSBlGjHMeUG9uEFTKROy/XorvU133zWVxfDZ3NkTxFluitM7
o8n92M3PyUh07slAR6HMyGjOH7DtFRnzkl5hAZ3d8sn+xiuGjOjx/JxJzNUIB+w7vT/IhfcEdwFq
yZC9Mq30M0OMFXndYR9FG/nw4nQnsYpboI8cE3ae163bUEEr4CVyNSGg+KwBKwRGhVO0JkfiVWYy
mzFA2G987XjJ3nDjryRlgl/JvJtUWO9vhjOvN0qh1AVivzaTWCwuA4gx/uzLIXMIi2J8F7xNEYP2
e/+UQpbZ5bo7KJPoshW7rLHgQz/zLwWtgnr7hds159JHJom6VEwOkxVde55RyT/h8dgYllz8DAUj
D9K3neJRizgnQFZcoAJhU0tuXGpMZHxu9dN/fv4qZ9Ok8DnBboqqpzZGjkk+suNCw96fCld28LgU
/yWb+bys5sDpNYqTXTceyAPKAK/zCEc0KKjO9WE7QW/WAMmgq3U2IJAeCbSwMuFALb/b7ahjwNaj
XVq34zh1oGgwRyjjJjofhbp0yIDonS/Qe+riW3PQFgNQEsrPZaC4XdzI3wjsUS37Z/AEnb7xys4f
5FIQva6NWIUOL849ArR3+73Tw4sfYvHYqZgXPZsb1dATl60/L1MYoQdy0l1zVUHvvnzjOCc0MvtH
l3Lu8HOQBifp6QAhrwvLzuGVCM6Si6Jh1Cy2yGM6iKX1Dk4BQijzcGJh0JQBy0O5AjF264Veffi4
XU7Tppulxw4GODvD/cPdzXlNebNiTVOfdDXhDas1Yq/MXwaWMGkTG/W4cxA6Nl0g9N+n/4aebOEM
3LvlrbQqw3pF54gK+wBzAus546T9qP10JrWJ0a8jpZ/SkgqYsyjP/l8oUQxeUxR+08WDB400BMhp
QAFs0BNmm7iCZ4ngfq3+vAnQo4XKfyj7e77bFeNk9f09JejzxRzWkR3AGUzoIkD2dl7g1g3clxkp
wPNGTkUKJf9+ZVqfZXBK8RPYKQA3FVW5gUM02yZhHkHro2Y85llVe679jKJFOINd3sP5Nlt42XhT
ohyfzzJamqZn0fhkiTUy6W7atKz630T7lFQ4V8WJ9ZluIoL0mfMTLnMSmjLm+KnCB18lxLpKiNyO
26ndNwFECsHdczdz2kIodL/XkttWU9BaPNqpdJHLJNw7MBx8j7qKGMfD7Do1wq7Q0Zmw8qNbwBEm
joJm/JXHatAtCkGRMn5fw/C/apoShmNi8vLSGZc4RnZvCRqI060QYUECrNtm7RYcoX2zV8g7a3Dj
YKyIa9DetMejkuxMxy0w2Irrsipdjp2/dqhlVr8laOTNvnuMS1/4r0AsABOlcoNNMLsaqm2uPEC/
t7ONeBmTNYYz0S5L5nCKP++eONH8kRAHRkeWqdasdzU5GTVe+wopfElg73NCX8BtmM+e0R4aAN5v
PTkH/usPSIe+7UGs7w9vZmAqSrUWJjD37MST1hDc3id1m2S/tSXJhTAUwLcNibqh5KWcK5IG2hH9
L/IvnNCj4x1VLwC4meWXa0H4KzIL2v0EwBruFNJXu3BCKgmL+SllkD0e3kfYQSILcHXI7VPCSMvW
11j3YNcELFH6ZRfWs609coYzzqdYdGkTL1qFfPZbTgopzmxc2QpwSjwOibnt3F2o+fiCIen4AQTK
45OiHk/0td8dx7xZqsFTaSAPuf5Vq0UUyKaZzXMr1fanhMd+Na5gjRbos2LMRZLS2Jxqa2qj9d3y
WVcIu5cYVc5Jg+INcCH2Oz9/uoWkD31Rba7KtfJyz7vH+kfaYFPKUWPGpO6Uu7hpgliLhNOjX9hh
fMTgx/Vo/nR2AT17mhPIgpkoUSdb5mtnw2IMF2q/KWi0UBSQgHQT6T6tbv4zmpxdxOD+dMPax64z
OBmC4ymckrhxOlL7Sj+vIRn/xfsSaOy5aKpSMrDLkiGYcFB46geStmJ0jCLPtxxBPDZQWPfQ8CSF
OAsu+A5XV5P4SoL4dHL7H/7lg1EBFTnw7wWzu3fMU0nRA7osjFQALAP0NWE73YES1QQ2aslvQ9YU
KBHlugZPcPUJX9s80TQqbJnLoZqR4OhKM+qX9NPmg55OJuMrsFGxdyktjOe+Ld24GbMIHNZwt7eA
1uXOq8TVgvH3o0ziGcGM4YJNZnS7GIPWwQb+IADX7wMaA6PySQONDUCTojdWn0BVeoc8CY7H8yaZ
yFqPwbWhzYCb80syKHFPl+4yAfna7yfGle1yG0SxEaA7FpWiI8DgoI7Y+7XxyHy8EhcXeUUSw+H2
88fwwOn6kzcQFvrjp7AD0/ennMYObDfaw2c00552qyy9H738QT/3Z2LHntGp36NDgR0PXmtLMfH3
aQbSjvOnmgES21//ofOeZxVtpQIT8Hv6ZqELcbNTd2Tucu3JFZPUMRWOsoimRqPXj8x9YNtfxNHm
70SGYscud31IxkjddmMrPsAJkzD4VSc+i/ri97b69l3YVH9CM6a70BDKgYJbNcPnyIOglmALgz9d
Y+7HTncuyWO0haUfqz7p3TrDj2q3IKtj29jsHXExBwIG59hQ5VUitaPZUpD1EnsytfKholWctUo6
VRBe/NHrLo8ELywtlmyciDm8vbe1RobLdIeqUnCzj1VsuzTBLc1oFbuR2VnFALHHFz6seve2H/sg
lUQDRdIAP13ENBccmOSpLbJKkFVvWlqY4dsMjF9RtftNGrwj4X5LZ2x+KQ2J9RDTAdhwEk4w2ow9
4n79T/f0ZWUUEfNZCTS1n7wA30CdTb5+5CNfoFFy+i2CC6SuRqZQyTjBV+CRwoBkIG81BR91AtIs
9Z8qKZGzibr/DMnXNxzmx7/Ab5yzM2I3ORBcyVoIH2/djt2tmZImCIxpEF8STaZ0rl6iM1lwJofa
pI0ivPHHQUTYCqZGsK/+isszt1KTTZzQFXn4KJLB6UADxZVebPKBnqIpCb+JhpKy4qWiNADkSvNq
PAIbSDS5DuEcAw1tfRHxMdd2sg/RgDfl+m35Wf6MockV02LZflmpCBAFO2GpyqAX6nEiuW8/VSsr
zNv5VBf4sNF7mwC0qanc3m31lN49qDor34LBapNYWDX5rSNV1JdiDRhxxeWcCMOAIs2qtMdL0d5B
WC6d5AORecqej3Wemzb/dWT9s7C+heOkvsZokLD+33EgJ/4tMOWE5K9aOO/7ZGuVAocLd4yNvyLZ
3lt7ynwV854tZ7lMmxgyh2ZOuEv3oAN+OJbD9H5ZJ5aAw/I7IHAfs7aqvYiUa4gxh/fQG6NJDIlO
YwI1AzqXeTbJyy62+AMg2voieC2+FbAFzF5C6VwAFFsXqy85Lo/hsmFus/aHpp43Sglyvh/cg4S5
R+ff7v9DMAqoP0TSRfU3JCyQ4sJjvO8lhjUOCJ56g2iUAV/nzUGF9ZVuKXuCmipDb7uvrxyuEr9N
eVg4FKG1xsuAraOG+RtZnT5rhWR9oE2ihmdD6Ync/rmNItioYQft7GsgoUVfXKmRlRqz7vu0eElO
a4S5fsKgPRhf7rqqn7URB4EZhfkXKx3tZcboMb1Hbi4p5K0orCabhpy3WhgLZeBo0b8Ag7ENyM7h
VjCxJbdtil11RXRGemUvyGjTDntF1yg6XMEE77jcFjNX5ltLcB1WxbNEqJCkTAGCBT92U23JCX5e
wdhHuxeIyArdPwQJZIyIbWacAUMJlR7LArX5X+G6IE+TQ50tAktX8Qf2TXftHpOBGDHH9R8KR1cm
PAjuU2eJabcBpwJPjIZN82m06WNSl51C7vQR1O7PvN0osozzABKxR7JyRFqJIIGPtkDxjcIQP2TM
qta6qess2vx24GQHFQKx2eLCAIVEc0yxIaPLvCzQ1krDPNuPzAs7vL6kAMUAfyZybvaOdGBxRVn1
RhJfpzQbWd7XWRLRqck3++BeQOXrJpuBL2C93LKDmuGLMqadA/xmgQZX4sUabDUlsBj75yjJW1Zz
R1K2baEy3AJyVdRGTV78slTXp6efFxqM61cwD/Sx+hv1p0mWqy2MlJw5ll8wIKCAEDYWfbTfs1cV
Qle89BNJQgKhJUeRStGUYrIGA/UZCFvcBPVx7LLN4iuBL3vEY7+OX02lvACYvOpM3GQMmWBLOLKR
4xVoqc9D01FfDoAO/TgBB7RtuMmhq13D0kItdWvJ11Wz9zD8AhPIA0KJ7QUpQsM0sCPEjygp08zn
KyxKAo7JpNIVu6bQ4yJ3CayYwuZfa5lOyCiIfwU+XecI/wF8zi6LuNudmtgDFzjxhxcaY+gqXRkC
MzVgsuk7l29ywXIFdatY9/O6V6FYlL9edAms0AF9VC7c55tqQi+iFoGin4E8Eh4hXhTFJSeZUSCS
goTSNJ89FW/pzTzzudXLlCN1j8775aMmD5yj0M+66a5TIlUs0uXmmDCi10eChQTV/LxxM/jbYy6z
N9Ve/6ii/tSHcZfAcOfM/j2kkaoNwWhKh4GDTRbnW5AC5WRFtfRNuEdbypf9pqWZNtZstHK5JXuK
LNPzfRVWDPcYXsb+/9lRpqzVhd6NgA6gXYgRU1vAL3a9FEXDWphUUG0TXWAycV+1c0UIy02ENEw7
01Z21OnDxFwQCR1rnswi5+ejVOqiFTiop2VTn49zdXShup7/l4Uwh52q7YvEjcNp2xUZ16Pd6tsJ
W+ZFPsCaTeRyS2bJ2uKZkKzHfjmmbTck20zBcD7nw0cRAEtptgNGroQ9tjMkOBVLTHzhCzeZZF6w
6VRHdlDvX5zsHmYzCC/cQX8u91ZoVuAsN+pE3WZQplZaazMeX/VIPP0WsDJ8cQGUDh9kw0Lb+hud
Ts9Q/ObnbvrwaA0CqQyvK1w3AxnepkoKBjZVJdAVTlLANjIFz15dBkMFHtlm3sUqurE7xlRwxpOa
DLGFXizOX5MNDKYmQHbNsn47/a92t++fcHn97wqkn8aqNmJdoeGSHBS/BiiXU8RvnnMnNbW4ZY5O
WHt0kTqttf0nC5YcHfYb2qy5oC3RrcAytjo9SgaIcwRhmYlqjeP2fpUYM+y9Oqqv+ilLvaOxEbka
UiKpVr7WJY1731g7LA92R4snO6FURBXsEur9WmNzrF/wJ0hFWAAYDF5tJ+uAymo8hcJgManHk3Ps
7lvUJCriH5XZrCXQgKlvs1ZPok+VivUPOGV+DG7+IQDIpfyERAINzP4SgxCb2/aBqfLgihR1R8MO
/eSUVPNj2aJ+NzsD8JHabBQfSSEKdzPUhwp2CB/XtfACpdPlM0wi/i/1ifTx/XyYI42Dghz4PG2b
kIPD5Di7fXnx+eaS/b+Dws0kBh477a8P5v7p7qeizlaiTN4rgLDHdXR+OnH8mA9y2jqjnHLdy/6Q
/FGcnxVY9+/lcEfaEjccZ58NP0JHkIzgIav6F2bfWFwlTw/7CLz6FxU7fgcpMruo7LrSWHNZtn3h
0BQGBQEucu4g2x8HrljnmuSKXK/+qCGwacQdDeEcjCsIJ1DQTrkqLX9rWbIH7SBSIOUPJC7R16eo
6A6OkkOkI7ZM4mJy+btV4GehyqqT6/SD60NVCIQ07pJ8FuzGPnc0PB0p1+xHvZdqFc6b6mfv1Phw
R8GDmrrg2G7BPA1tf5q7rmZwULAkpStTguxaqhxAnI0vxGkgeBYnFC9LRKDzRbUgpZVTrsSqXMOk
qpHycXYrZMsJDnwAktWaG4E9qyD3TVH9vcrwDU//TmK/ujkjYWd0zPEX9qXj79V8lvP68AzHfYy2
YRSbgi0KfA8tMZWzZ3iO/wevgcI7dzDz+DqqkuCix5St/+5FbyComjgHa/9k69aDvgd4bhCN1YOD
9EWg2+HA83Zpk6cRrfyS+yZrxaCGMEeBBao3dWq3gpxQb70VzyY4Zidf7SJOfXzgvNjlnYfOMs79
r0KebCqZimHGtJCAsCKzH2mkr0hWRrAANk4Lic9E+R2Tgl7KQTnAxt5b+HDsyp5LOr6d9VKNV+/4
nOEyzAUWo4DYQp/MCdZY0ctQdmHvqGFhhzSX5BXRYoh/itnKE6mL2Zt9ofLmaoxIGBh9sdH3mx8r
2RS6VoH/mXleTduy86qmgihSFvAnKbvl96vbY2QMHIn5LhZ14LgGpsI+1T1RFsFZfatWepboydys
N2vcYkE7MU6z1/ogRXThRneGlae6O/nnLnmWQ1AYHJPb4ElkXQTABQ5/jC5kQMAAxo10+VY3nDR9
ntDHsY6q5HSVZYIDM5dpX2lSh/cKD6iCYVU6y21eAQFnHjkUb4FPoAZxIg8cpkycAsW5dXSTsdJT
msli9Y6EQQKNFlj5gNpXDxvTq6isxznG2LtwARKrv6h5fMhdn2tfufEBTdnkswFl7iXODJdYo9xT
G5Qva/LTa7qViH96ybzDlp5M9mfObumr2CxTOU77nL+SJHXCg+wIDbc8jIn8nqXUnx8uSUfi/kXG
sTtm2D3yHxSbks+pfB5l1Lw/ARKa1twJGbQP7/uK6q+I63KlIGXgUaPL5IjP23pzVgFufEsue36X
m01cZgAZciZmrWvlNNSU3GdfWOrOkXdZVkNwnsQ2qd88EN0GT7zUI2lO0855ryUC1LAxhRkr70qT
8KfUtq2aRZYSZzu6PNg//UyP3YSvi2ho/eQqJRp2RsQZ9gzJq94NYapnPBqVbSmhA97UFSGFmBI1
uaS0rfFpLplfoJxs+pjwk/ogKZRN/+7HdtXVlf4Kg42iN3myZUCIXTgpay+PCpJaGEyFfBFhLE2d
HQRd2lWZsjnyvuAwOuTXkE5iiAlmRKREBGbAFiqVR5VgHxdwLq0h4EJl9Ascrta5OwlulnCf6uMI
o6GJ8uDWyQBMHuOV5/2T85/V2F63Rv7eqTI1WXEAcRQYSmvMqWFgL+t6dMkriw9uhUtGe3SU4C5L
M2gKwgoxIrsUQlxpXg+KMfzK+kdg4zGQuOZ60664q3CHi/lfTZcFA2K5xwtbhck0WeKwrvptJHx+
GVCSxBnws5CPOjZfvsFGXBYpuBWB5bbJcR2dPWpfhRqFKAQh1BVz6xOImqxAeR08FYV9V/eekMVX
/8p8C1w0a0DtiHrvpBUQJ53vcbKqtTTvfniiN+OICJX6zDJmJlwUHeiGbbvy+uh1HGXjY4kGfwO6
sSY1SVg2iJp4XATOuUxD9AIUizSkPtnpsZzu9B00ok3Be28v1fLVCz/hPjdR+JT3b8WnZ6R+Ue6A
fxniEWFtIi5iL3egBn6Ct505NF0SzPeDb7XGOnubaGRJWPfMUfZKRwA4mwtl6YTvUlGR5qkNSLby
0oynbo/K543U8V6ij5Iaamm34VraHuxBAVRLsQlwtQ+yoACBAeVtkZz9cGVBFyXsGpDO/OPnN3E1
2SIZjMSGRPgSMIYcSaGBT6N3390lPINV61Ocfm2qZwuaXCQ3C0PJ6YneMOSkYed+qgCr8eMMmVTI
zwr0gMnR8ymlUMFG0OdW7laAi7zwH/78HAWybgL5TbDkZXUBMqBHixSCxRSt6h0/Yiu4a5QTmzwW
V2wG48z2ILYdcAO85mUMMbm77itdY9BUGfB3ZvpuqS8BA1cHsMl0X3Nwr7SG5yIctKv9O9THE8sV
+Jm2sF6qFLRuS0E/AtLLl7sUOcK0w5yNU332S75bbiVSUye+9gzuMzMbAIX+UjW7ckQNjoWHsXhn
D544HLuSPX5HdSbu5Evb+2VaXCdz2UnRjOd2ZTCcHOSZfCwTw9bMvo25K6oRK2ghHXyKKB5UZKQK
6L67DQJHP2GNwDL6hwUTgYpP3Ta0pwITXJBe4O92y5JTtLKGb59drpUp376WO5jPSkXP1bSx4363
TdBqxHOFx7RIiy+dcUmFgAZ87hGHBuicQkJrMz3mK2Iue+egp+/W+KUZqrKeJ+aKaGAyD241OmHA
k5IYjNGqfqW2FKwqHBLQUSViWOs/3zFWdawITymWbXs9oIziK27R4nuBAJxshy+PsJ5AhGdCQeEs
CiZvmQcmUxfs/iEn6iKR4mciLuA0jMAb9Zn3zjWG+QGGOj2KmCtm6wXPj+ryUK5iNXFhn8+6jOSy
W+R+2t6P56FTRtFmfUktwgHA7jjUTr58LJjXjSGSIXQsN31kNM1Tl8w4oR2rGl7deWQE+UUzynaF
k4ebUXvwMOu+/j5wT/oLjw/NlGlAfmioc7FrQsQrf5ARv85gmKBW9Z0As9xFzjbOvJRJu/EPALFe
7+Ccm0HRSo8lyJSKplCsLUCt+ZW0Z0B3oDLu78ukM5bdPbi3M9L1LA0r9LBvZ17XX1bDrO/63p9e
RxnxAEinkqLQAGNcpVwEdgohSADB5I8OAe3ps0FW95D8Ln23dWE3f08thYLZZhy9hywdlCbo8uzp
RwIsOcucwjCHz8gn7mHZw9f23/URETJhq486m80u0OYeKgV7ny5jZT+/8kpQWGYEH8qVwYzFGlzZ
b/yJX0qZpD10+u88LoBusm15k2cg0cKgPzhgdahCBLyzmuHx/bkVSJ5wTj2rIcMHTluEcsdiVIAw
JKcwCjwiFdeX+iicG5ocDBTDEU2MKRBH8G/j07iKFEcyl1R/9eynLypnCnFaYLqZHeCcbF05SaFP
Oyo1ZeeKHdvs2rkDG8vWmVkraXuahcBy+IaODgAVOgKJ1cCusHdRyRBv9oE0WbhDvIFBOZu3t311
bO1ne5/QhdovLuHWiqJ+r58vU3g7MfcKaHTf/BuP/fCsdLRXRa34Gc4yDDjIOB09dhWRg2kCfMTW
jLR3z+f8FbfvOzRNBGHrE/TI1UKsuQN72MlFcNbMV5Zx5ALFF04q6mdzlyR/BFN5zpxuTTdRUiXs
3RI8K1xDP+6iMIS9pYPfcYLFA1vkdoCSCDU0OPfKFn0gu4ctV+jjAERGNF/527PaQk/D57tv4h7z
WHwvMBSxokUUJVFhLK/4YyLKJqFDThpZ2HAkayDzIlU89FCh9VKX5hl4zweNINJhRV/yCSvJDpe5
JE2s1CAav23p1rLimSTcYku1AWo21oE+HK7XPtfmk/npuQvXRU9xMf7cfXTYawtunz7qNGKv8KxJ
mK5OyGThTWjkWB1XZE3/T38sb2Wkgt0xBXvqsUT4egl6TbJ5e+RiLA1YHg9mbv2hdiMtFJewxoMn
6e1h1MRVJZ8uPuZHYrxZX6J8abCobsBCvSeQ8dH4Daoj35sg4CLJL5DYBCmqo4z4jCEbxiruIQQa
SLeVe1OWyKnOZfsb6WvAsFNJXgulIlRlT58BGZm0gqZ3cND7iw9367rRMUkCvoyi0dxlEvGqqpxD
uIuqQP/sUp/Lz3Mz6Ct/MzfBkYfrwK8/HXfPaFLwFkPbZqTk0brfwEC9YEVxI5Uw6bIjEkWWaQwL
MifFosWtysxMHKOtclZsD6h1RmrGmoo9+szbHIzKv6hjzvxtm9mGqG1r6OXx6CgL5X+4Gknk8pvv
zRyMVcoUQapboptXPKPFpwJL2ZfW5F/6lPxY4VhhIRGnIdRaFrXSjaziLaZGATZ7QAdUI0ZpTf4A
9i48YyVOu+BSImlro7T5uuXNqY+DlmOxqbMTDRMr+88kHmt9wdL1a2se/ttFVRhTitqKSlhfXSDM
nyK/H8asN5d/5avlMu4EEiKgjsVNq1yMjRL5AUoa08fsGjY4rUZog4mhidnzb0We3HaNfLUJzEsx
DzPFWWO7uoi58Hi7Ab7j9iAwgc9rq0GqQ2llSloIpyNnm0tcutcVFwQ17/0+ufvlNRRk/R6si/Px
MgOur7vVjr6cg3Efk08t1V6EXo7KAXs/qjf4pkXpsuc/4HVoinHDMscJcshvgYAQP697XmZlx6s1
q8vVnPSZPzYqKHPJZ/REmgXsgNJ+qrNkNZWbJzcShWgDTaphZqLelctzaPkLuiS9AE5rW9xP59Ea
Qk0GJHK2DpDdzbXAHHcMjyKinq9hnApe9afScHroks4FevGfd6QNITQWpoS7hWyrDuIOEvFJVMHr
cuF5+NllWE90KIBs33x6Vm5Hp8/fYkwqzLoleZ8eqtEDe2qpoCqYJXiI1VosIZj+qnpITlzthj97
BDGdQyNxhlhWVFmdS+Kdq5GJmd7v8EEgshv+rpFjjvPgQlV5cEzvKiprVLWFLLrfARYS2hanJ395
Cnz2E5fp2mvaKo8G/fLqhfv29SEGVpLPRP0dimQEDkRjllkF8MeVlVnwJf2G5LkdqHAc2tNhNX+O
zC4CHujUwJ5loYvTapAMTXpstPoWCcPk4vWHKapgVEy9TynoAKRZeiY/NDVdo8WT5WFxqc0+Z7t2
hqsel3QbIvOiHcL7P7P3Xj0LZHVHWzXPHtWI7hwad0OThGyuOKweL9hvQajtRy2hLf0xTD+LaivU
j9vZQl5ENKVzvVblAqJ5c4gp/mmVaPzev8zcSWa+ol//2mHJBtK5AzXQeVd/yuIdsilwente9AFt
aQsl0VHKwBCLhnXMaM6L4l9SJqV7AepADASR9dbZPKRfSMl0loO3kVJLXBNmX7+u8vK4GJEBlhPl
M8SZ7IEvKBKNr4NxQcrYk+qgcNaHM3EULXgtpGh6Jv8+jgXS66O2NHHEDyaR+aQYPolXcbxFl2GF
`protect end_protected
