// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 14:24:35 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bvKa2JJnFFXQvFqSu/yMSTrjvcKUU/bFMkvFefoLYkgEtBlv70dFRad+ahBP5ql2
CaCQxNItKZ8xoVKQgzBQh9BLZxw0HpohlhxqWy4rpGEZFDALlI+/d3P3jFkqq7tL
SIAg85WHNyl74M9Qq9ru1Eq/01Jb4C2mQuHk2SyG+z8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11200)
b4g6SOa2jM77e9uX3mOT2jK5JCZeUgrm9bQhyugJvBUD++LzHMKBn+KdMZwZ/I10
DrQ6QNFZ21Vv4/I2AuVnsR2H5SqiWXaOgYncJHdt+oxzotvvnPmYh7qFrNOOPwrk
iebS7h7yaFcrNlxwt5jRFlL6wEAR0nZXgeoXI+hCd9MtwV01ALa9KGotXpTPzgFZ
+6vi+I/zqP/jtnPVqPHLQ6s0Av24kYL9v7i3Eg3hyM1cQS56XkCOqnakELDcMLWz
PhXZ3PKL9RbtVAHnQz+BkU/ikVfvAMepfDzcJLHYLvedAbb1u0zI25gyOCrMWT4p
6G8oT6+gHhBowbblgUanlGB33zc7URlDWavnKehk8mysHZ/P5U3UWE+B0ZrTEVeN
i5xAUK429b5JNmFxYj/QVgwL6hlZJExcUaXKUUthXstK5R9Si4D3p+CZlQq/skc7
uNIBZDZt5lw+xrHn4LWH8iwK8+7wb0GMMIcvHs4QH9oWF6XhB9nNdXkWz3tF/vov
O46t7K94g1lNZJxZn1bJvTGdod9ZcBYYZWSIZLC3RaWpEMzg2VSdW0DXgVxhvh/a
CpnobnOjnxQP/chgsKyHvxk80VLW9oHLrkHAx6g6eRKf4VFvF3NiA8U+s1eUegG2
1mOpXkFTW5lj7DhXjCD6pkwpBy4gBoWBeNripIrSMwSzzppMVEhkPSkY3zLWl7wm
YY+gNpLcrnxu+aUdjLtk6gCjFBi8CRl9jwYjt/t8NWHYUZpRBxJe1rNq7vo5auEb
7DH3evuZQMwRyDb5PrFNBXpQdKVNy7UUhm1IT7wGP8QXC5Cg8FNfqZw22kMgosCV
JdmBOM6At7JRuIMT/OimuzMe6jUBmhQJt6sH8SY9IjMO4QDSBqrhN75WTCvDO5xx
DzYePQ61vFbTowg8k78Tw/K68UMiFytiXNSiROE6p0bqQ0eNRaWmlyKhG65ql1gt
gfOw0+8SoqioElxiMsWKfa01aD1GWwHzbYgUtBSL8ktwg2WUzxVD4fgN1W1eF/Sx
oshN6DVhzroSNNkYwC+6TIicB10BSBOvLDJhN2MX+YAfbHSI7cI0GmTUpnZlVlcm
8vJwLs9Q4ywJKGJ5ytayl3HGUNPT/xujq8qUOeEI8q3isaDfEPaXfdyvCT3UVl2S
RH4jbkIuZpgl5U/iCtpcPOYtBqLimpKI+8ClgdiTpVxAYtn4Dq4Qc0nUIV1ozqbJ
41+ZG5JXlFPJ32ZL9E7zEI/ic8T1uD0WqyP3bMoQ4AbPOeb50WEoXv7/PvV8KMsx
FL5FGm39phQ4eTryHWG0oueWGavTEIN3wxUcfy6c5PUpVDVKvS7j9BBpRKJov0h9
TJS72HuabmwQViLWvHDjSj6kO3nHCzWpXYi0VxClIf3Yvj+g5ZpyDlqMWFfl8xJY
nhMWLrqsmPLEWmh62+TgxS7wtnDEl7txqP/MAPRxFiKlZjLXYNWyyQdHuB/QzHj8
CHx+bsE7Vae/61/YewoVkgll1Wr0QH4FfY6cBS5+s6ej9U4da2rg3gGMLeFloMe8
Q2bE7S9FfiT8aTYq/viGRQs0jSOzZbHQ0umEvBkmOOLAMnj1Msd5H3vSETfR2IYi
zGRtRaZv66w23j7S2tMVPDqfZba3U01sgmWjzTY3qRCKy2CiLE0DDm3VdeZ2j6Vf
baQny/3kky99eojc3dcyJV74i9ndiDF2Cw8D2x049feIHrz4otKsIT0VSTQMzHqY
bMNuvUowV3YBnCAy5kdUTippp5Cz7O1SiMnj4aYJPyBVzt86POvfoUD31K4yiVd1
enJwb9PA7RE+5JvEBgTvsjbjDjgiV7MdA689lfyxfaoQNgrS9LutII8DqRWaZQqY
+OjS/+Sxgq4U+a80EdS1AaAwtm8D5LGLNiXif0aG/my0GPI+/kKybhSl/Z1ydRSh
Wn+6dDXJzzs/rDCjmguvEwwKayo24tABXm82G5L8PzZ8XoFnZuTvLeR36H0ji6FO
LeLEyiArWUhcGM2kGjd06Zrz5FED2MyzgOIfO4ZVP3niN/EScR/jwqeOBnorv4lX
VhfeMGvC2GL+uEQM2oN3uf/ZKyt1a/WGxHKjyBgwGOzWBcCv7gUM9K1phxxGX/v/
ks6mUEdS4xJPsmjLckM3tYjiUaBo9z+EDwtogR7otyHqY1E5VCEjWan4V5hbDp8I
X+AEbgKsRkr/zm2xjKHOcDGc/DUIZ3riJMcgmS2CmofNwpNsRmw4UUiajQqEL29H
h13srTDDjBO6ops8MG6k8gSBNyNzWLsdJojWsyM7wDIjbttXKPdQkfMZepN8xMz9
iS7lqNaIof2hNbodraFFcLnzekE9OzOrKuonVX3+St9J7gg5uHvWfRAAR5kcjybc
BlmCRwrqM2zjd3d3FHRj6CR3DPgOdGWSiN5tcXMB8yWv4/NkGrsSW2vG/uERQiT/
3mCjc4B56EdHs+jyKAbzEZNZI/I7TArAHYR8Ohqi3s85GWjN9+e7zjUMZVG/RUa1
F21qo8m95LFBucHPDX9dw7em8r5LNmWO0Mjpyu+uZHVIQwTRSAvgpWWg3oifnqKq
ibHCCg+03I/mXeXO1Pb+fJ464/Wf0BTzlyZmkrNSAi952Qnq7DDv8O8wQOpmknlV
cQhTHsO1/Z45CHuluEzlnYRt7TJi24o43lwtUqUeLvLPtx9cyFyJA7ZSDtjn/eWu
IlxdbYehkPdWs8nid+BnTY7FlodUr3cw8VdzHHjgvWkOVb98nvMIjJmX3J4BIjN1
t0u9JqN+NRpKIgkw2lmRSLxxbovFkxL7XCYc7KQqB09KsxeAYCZIXvEL2pRPAhQa
5Cfnd7FdW6Z8tg2f5Om11mN5vFY8qsFNsDKuQANeqdhRyTs8NWniREI5RLEQzxOe
pjWvq3Fb0vRi8CB2fP6YedT2vYAz8NFbYY/8x7fuFkuyQOVKa72tqRkzDJduZ3d4
nLhpmFGMU5cHaarGNg5+hyfxJ6evioCdDcngXS9OpuaWiiL0mvjn08+7sNSwb6jI
ZHl/R1nlLnmBawXAbcXknUn2Wn1J6edN1KWfzF3CYIA5RrcDNp2WbHED/EjQ974F
GMfOjc0NKInTjPWA+1BKWI7ZrghYVItnZx2BTxGdwYRioy7hWxek980BTQjQQ2qm
d2VIERpYuC53ZRmceEH6PYulty9izo4dlGIXmsI/8vPGSdeDhWBbxeYubIfKbS2f
t5P5f+YapLrWhQKGCCZxonCDTuIVh3IH0zX6OtGqW4QG+7drDL2W+jzgViQgEdJX
jwsL1+kL/gJM188N6h12G172zyeHklDBAhx15VYWA4Jx2nXEzqnnjDjFbTPX560d
xb0sho8AbdJOVEkQ0dLfcNS1DE3G85UB2G64DPB74UHa5qvHYTogUeGYh9cnlfvU
EuXJAJUmV2R2l2X2Zjn/pPMnty7bUqf7kTp5dFmNCiRTUL1XKZupsfyTCMa9/GXu
H8pkpCrw2JT8Tcg/84RDkV7gmL5R5dvtC/3AGQ4K8BXK/mrGgcOg3lQh+r/DU3iA
tLQJhmzCfRXa7/77vfvnBLDNnoDaTaJ37eP4rGZspyLsTwxS4jUKC/MGh7vQSS/l
ii3PAFHKNOJFM5gEv6hz4rJrkiVVArkJ8XupcKNmR3x1hPVyTIEuFuX5DZGSCzzH
Yz2B430VHs3+XL05rkiuEruRnf1iuzHGkRiqvlMcwo9UWsCaVHDWwj4hpzkEJU3m
jwi+NrgdfTdkjgkyZlmH7c0n8ZMTM3OTuL7NwDJY+k7YwrKF3pErLK3rAkBoHrgS
IuNqt0fKIFkTSLMxCL7+VW+xMgW2ne6azU54q3auW4Xtpa7l4pBLrkkTs4J/IFtZ
3GNciVyj7A5h/UoLMjTpSUXjDSu6gpR+yrHh+8Zmb2ZzP9pe/EW13Suhp1eYSLzd
UfKYldAN0Wk7Vx5HQcxx3jDABFKt9yLLicMhocyjPZvuGHs1cIgbLNAJMr8iGT8h
jQi4fV6PTGcrL8VZtVmxEztYv8517GRkVaE1fH0UY02znw+9v4wR6XxdqL4sEqYk
WaynmN5ieEi0aSqRMauJBVJg1DDWODOucvymJJfvU9Fd3Q0ExrY98yUTxXzrFBwK
If8CHKac4jEGRZ2vQg2FWNlvzXlmaA0qdHQZ1Ea+cDouZTqz8mu5FeTQ+Nwjl/OI
pxhkcP0yndq/JAWnKxfljWrD1WysHH/sfgg3Lkn5pcYO64sL4JYaTIsfs4G6BpoJ
9dujUdmi+YL6c+TEbLQDi0X0+yO42ZKx8c7qIVGyVqknth/M+kBW92cyhFL49QiL
H8xWbjUgb1DmWhTtMgfqqjv3jZXRF/unsxy7jcB9CdO5IlUPXIU0n28hM5kto2i1
pl5N0p/NMBX/QmvaS2ULbdtDULY+x9gr2ezhvj/nF+8Tb5we/RFxvmkXR4iS+Tts
DnsiKa/IBIkUG/o46x/HRuT5LKXQCu+S2Ope53XQgagcK/2xYIY9g/drwqmjEBus
CLlNS9eTCYqSpy9Snsy1Tu5v3iB/fNavMfFLcwGKUqS3+pFRTwo4b4u2Fq097H9n
6AOH/YReaDj+kK9cyntIZGI0f5NLV9vDgKo6ugRnMbDumLtha96RQRbojjW17nWh
m/68/rdNNg5mUYgKQuqPmLDyZBswzJAxhO8hRi7FrDnAy+tk9WZ10SAKw9S33+Hg
MNOCoygD5k01SHYWVPVukyJXh227CELaCvrqtMy0BZhsm9q7tj/0y73slCIK5wa4
iqlqrPNQNcB7S4md0DayyhQUPETwvYVlu5gkvFTLeNc95qa8QXrMoqiwFo7SapCC
2A8kfraXE9IFrO1fDzBDqq7EbvpMt5VQ9nr/A7sYxLhbSSTWollUesIQH4jgGfzD
WXQBgXyHgkfdEpZgOw0TGRIhIT6mnvzneKr4HV45m8SDhDnEXYJj++6n2Hp+Xo/C
F+JhRco5NZUERAvDVXeHH5pel0dWZkEvaADo8FYftR0swy0ekidyp/dwVg70Gu+H
rHf+52SgvFxtM4gpAhVGtBUowD8XMlC/NOXjzUb5+vPWKYhe7W+wL1OgciHuvVbR
hhMYr/S81QMmIxn56nF6MwNGOh8CFuABkAJTCHbqy7V4lqkbMgpmWHPjcBHbJ5Fs
ZSH72aGQXxrCI4ZE+CMib4Kck4wwDZYD2Ht6a1l9b5GcvdcxOzc6rZjv5nbedC/C
bVUNQeXxGIws1oGVOkeS0TSosniL48snXW1Kp7gDcRfIiiGjAE3qI5+wz8O500xj
VXgLWpi0aqoIZbpjiPVWpCWq7ezFumBZWDVBq6soqCPSMGOufG2WKAoyXyYUotmA
wN+0rFOEAXlRd23NQy0HcWOQMwAScL2wgoQov2oJlVRHMHLQhNyCCpOlcGUidbWc
hCJW9vaLD5JlXjcJM7ipLJMpbXH+gWfbjVhB5UUZ1kyUNlO+5YeDXuB5KTTNaL6b
Xfv9VayCpaZcyThitt9F67dp0m7+5uNj0ds+77kRhTWsGxaubCWnvlaMYRoMim5s
KcZYXFyGz4BqHN2BqS2AFnqviO4DYU5YlEh8ZFalP/5ItrskVmXZxnDAnvNkIl8m
YLVfezSGW3NiRs6/C6/0dCzVGyiWvNL9BWMtJNeEZBQB2WlWfU4AsFRXyFq0K32o
ahijkrub9Ez87yQrnR/Ogbrgm0zEEeDsTJ7KonEJ+jchBN5+ZjjYMRI7r21Fmomm
kYf/HyPtmfOx6iQoP6mVrntcWpay3KHXyTHdbE7krhCa230igI2yiPwlqZon60ZC
mq5OOeixW8iTsybOmCmAtvc1WbesPcW91Pb87lrrU2U9nmbq1FhMzZAM+VF2iY9M
5otZSsImGqVxy85lTekE5MeKajFB8qyZiD23hEz/3+6R0ZzYUPvajiO/abj/stva
2Lt12weXAGp4LfQ4Zv6dUzGgeu0CEmZ6ByyTxjgAkUFme2npuRXeXz5FbDxca26j
MKeMrRIHrHUrxCcCAbuoXfbuToN3GR7oDsQfQX7IDRCx2VhEF1JvrFzmj4YrD3wh
LlTvFGFZjV5ZoEEkXwlydBQvnBcPq08m2JiHbfQiBMCHfeg00bRnjtcnJS3uPjz0
Nd+hdc4Krmbu9HKwf85qG1EIGFiK+lPaOFeC4xOVAJ6MusZSm89BuLyRXQVEJMTQ
sLx74rR2ZGE1M3idO0sEmCDJaTVp6XxWDivlknS0eEbBfIi4o8tMglQjoOug4ug3
MpPnuhOorTS5nlVnrMSVJQ57sCSZKmIa9OPVJvSNRZHD7mFlWS3kxD/ptq3z0v/V
ODM16+NPf36VOPqLFGBgbz9JWa/FPas1JJTDIBpx5bUvterWIVNMc69vyK8ayGxE
OOkerGZmm7q45KX5YQugMwYi3C68yV5Lch6CmMiFca0lCTsI2ONFenxDgN0a7DS7
HIacSuuB1qXnSmDqcBLdP9kNWcsxR7H311uLUOGGGNx79fU6fDSmn80JSgpPVc9F
9eBRN5ZS2xL16ytyLc6dxeLEEZ7PRxPCMxyQrRVA2TX57Ym7mfDbrr6MkSdkV8bU
s5pYrZXlSh4Z7MmnesbiZQ/+g692Qt4TTqVsK2+xoSx4X7hdtatFy4PI4oL4kYMX
4gHWwRg85k4z7oMXt0qbpvRTae/oWz9kt5y5jlH8N8Uph7v8O4g+EiKSfLpoJkcx
3IdW9pixjGWFtzMr3eF35RuV83BfwOEavBkwANt9lbQ3Bfev7Osn2xn00eeYYZ9v
5e3YUgwC9D/XsOON9Fsj4ZngZA+wMcSgf1MO5WmAJLUcYKFSR/wx+69kGqiIb0K+
UA/Lt6OURoIhnhKMT9EgjNLueIBP29ytJubBdRvgG4anv95cZkCnb1szt1wT/Grg
SYWYSFthQy/QGNp0JEz7B+yIc8LRuFvvgsG+0JXmAje1HIK7GRDQeUG+cf9NVJ2n
m6mJ/Go2wHmeIdohoxGJY7/5+SJNXVyWs8MG258CZL0k1w8Aao4F0+yn++VSIxlS
MjFfuV3fzqb7c6TD4aVr4Zsx20clX6qDB/HfOG1yc78w0pXxQ/leGNrSUVFU5+4l
5x/kBt6zxfkxqJaTzSg5bXyllhzTHrPVzMH+bOuO1KtoDySFWA4rO8o8mOldpI6T
zSViRPUTPKIg5DrQX8ydBE9Lvuv9lJWXRUbaWRbk3ALP/8/FJkPclbCggCrDSzNN
YK6BIBTnik1mEMn+HPNkRHvUS8/oKuYtAFlDd5UcwrZSIZAm3mWNVyzZo446UhUd
QsMqday2Frh3VGG8PCuGrm1sPC+HfJ3eGiqsCwsee3oD/uRaMOHB0ErKBWMq8pLp
JYxqF1MNMLx8PKL062v95XRAUBIOVwTtzmIjtoySqoGlsRTbxawdwGW7Lx5vEoLa
gcszyMXsSi0Hw2ER/UmwEZu28QmgkUCX1rHf0wk2iBwmMjUZeZJq1bCKErhuel+x
CNYy+7B/HMtLVQc90GpbyeCFl49VGc3Es9iZSw8Dn9Ir5ggtMikxt+DgO3JVGOHo
4yLSfK/4viD7ThcUxofkQo4ZNMEJp1a6+yt46LrESx53mACF0htmo2ERmAbnLw2d
OybkbV2sq2Zt3qigV1gOi0U9ftlb1EyF5sZXBA50Uk6cJX97fmmLwoPWHye1jKV7
qXCPQ03DBRUNir/erzG5TehjwGA5ibuEGNqhvNfvgUcxMN/XeCJrvT+sYU8gqqFC
dVT7BynZjzsjenfDQDtApWaRLCUvudBHP16WeHvmZIlJ2KDqvItgx4yhCSRmA8PG
+yWVE5Bc3G/aAcWLoSs5CKO99vmXfcvNQSHOLqO+0nvLVFHjXcbiPcUGdlacaDL+
U2CXI7nl98rPd0cIBc0n9odltyyrM7R/thMayCteMrNy2bqH/ak7f983O0KA+kD1
Klye1T7gmG49PkecuXMUnHQZphWflwEHg4dVDPypoj63Jh0d6+vuYjSgpu0jlyJd
SGDqgz3+RnpO90mZm/AkpRzwHEJE8qXfHRcQsEzcCUkp4wM6VQBTpKzbIk4DyMlP
qJ2Fq8I0QBh803ayfO6Bgs5B23xj6xppikmgPpBMCmtin3iTYcXwoUKqNvIw/KIv
B1NRv5Sl0s3KRmFhzvvLMvO51S9Du0cMliLfn9kCT0J1dn8dkKbxo2zjKeUVAdYt
a4cBicAqY5nzlW8w/dRCEylLTLPUsOyb21tbjZmBjge32zvUDqPwKJt6A83Kkf9r
5f4SXb3cX3v3Iwox1IfsLjBoqEkVXXfS105280xQ/+iymp07rMUAc3weT+lSN3Lv
ItdgzeJPYLNqXLlwaHko5Q1x/Oveq9J/Jxfq3paAn/flqkPasXJ/QKPbJZu6A3BI
LECP8xDTwzOVOjGA0oFZ/S+AWpqKXOlozqm3AkbiX9vbDCINsGVhnWPngVV3DmOX
A0V5/ebziu1AzJ1SICusBgScrxYy+VEuZh2J2NckooxZ3uQMgcKwOC+V3Ko5HLNm
iEujUp8v5y3WUBSQcOBx1BnIegV5b4nTv96IbZ24lPKSNruZMeyrFsAPh893WDQK
DYtAE5So2OtkXfh7xjUKLyANaPPjlOlxQnIuqvgtb8GX2lQzdcFL/d6mA75ksYdu
yB/mKv8dIeWltEfhJOgmtm8lr749CH6whupmHYlOfqWERnOG98OtBHa3MMQBNyab
VxPG/YfX6CbSl6ZEQ0zIxFcwPy8dJTO2nZJjSOSUX4pDZ8LX55kgS5wN8uFU8qsU
f2VKTU/zVluJpR3Nqt1XA32/L28roThbkTGZfEvXuNae6+t0j7p1xSpOrFyGn6qs
UAVivbScsfEZMDzuokQPZw/9RMJq2gGQsD/9RgtarDa1nReWaUweUtXPDeG4PpSF
eKb2La9NVJVFG7hEWkHb/8dFMkNsO9zX0mKzFKbEojVqTFfPFBovYMHVUgUo4Xs/
wCvpZt++C7JOJl/uG4HkMxye183weXu/3T72LnSR4ne8dvzLIEp9cBNvPBQcQgPO
UJpecxgBcAp6y1dkNEt5F6qnR9jG/koEQKKvzIQAjXRDqv4sd4bff01b8tuPKGDS
YWhPbEiVmASwLTJoZCAi/hCW3aJUyhG7f/HAgCyaMraaTDdYl8cQiRp1BvwXS1N6
v1lsG9d8ZeOW1BIfKE3JAS1O/0pZLt9jFNUtHNKDaEBH0E86LjYeqxytmZfNyeS/
CS9N+ENKpmuiJpz16mH4+NbRi19ye+3jSdPo9mYcCXKf0YNdn2TCqwLAU9KWssJz
wtLyGw5XB6nVGiwCUI7JblM8DEBja4RfBiLaLhBUI9DYc4mNoAYasLHtiFHNaJiR
Q1rXa5x6UDs5kSLOtcq4HLq+TA/pECosCP/N1s6i2E07p8Kh5Y8QoLyx8jUwdFkZ
duTUrVo+Ifu1aIPSXHu4LaP0ARqjC3zPL91Z33+BieFr7GtD4tqJ/bnWzpC6SuMd
91lwuFmXqQv8Kt91XWw/m9MNY3Davt8kyaWR8DQPlsiJy4jMChyxA15GX16WUlFN
NIVPn7g0LnUt4mGHttOhmLLYdJLwClOsG+Y+rFhQX2Fyak1gRE6IVFCXAyz/9/CN
CvfEAJFGxPKEU7neUZhecL2n2JShAeIHvKO3fuGAwUWAsnCSWuKbKIq4QCLYA5EZ
TeDKHMjO90jiUQUW34btbB0fEMneRJJ98o72sgEKRN8ko006wGrSJzi9Y2lV8L7y
VVfG/2u3fBglL5DAT+U06DiHvdznLEX3WlGH/YAkZtKevH6hbCmK1PxYzGXlgn7r
7jlSwgB+ZfhFiUBAgT0sVfQB8zJSSzMZ9KBDLsY2h5PiGR/S2Qiwdl3NCwu0Kdg2
/UMgcQkYfaAb4Lb5TXp9fOnWyzyIqWcdffsRmu3LxZhc06EpjN4+q4EBMAg2hBUc
IyowYqC26W9cUcJuXxUqQ39hDHGzX/A+701ydiquhLk0LqThhPN/caPEFNBGuWwG
mZAlytb1yw56ph8dUD65eAaovAM6Ps3hWMFE/e9biqQf2B8I4Jn0p96HAaYtmxRs
ds/LZrWtRkQtPme1787Jzsx0LNbrscQE2Q9jskG+T0ByM+rc/nKffNgBxYnMQv3I
+uocOfg4ZM3zO2cwZfcOaypwcT61dq7sRZ8pDlLGz7njQ4ovJ8W3+xQWHcbaqZnW
PJDrxPXHunaZ6FD1IRAtDSt17gkOUZJXK9uJkY11uOXXPgASh1YBwXjMcb6wlPmc
cvQSjIvqPZbPNA1+HhmFfrKr0uMBDATgzLuRNyqe+G0y2AyehwF0YJA7s0ivLG9s
FW9T6IMPUPnOL75mFB7UNFUgqTxFljEf44l6OI2sg/nWFSuWF5MQc5JJppf6Z3TI
8kay7gi4BxrpUdkRqeGj6iXLJXTLljCBI/1wfIRAeloW4Y4aXHtc35egWM7MxsWE
Ney8daL7Nmdv/IiddvqdQzXYaVTRXTMKJLRzA8KQOJkm8LwC9C0NZ7e4tR+1xLgT
yoRhkHFaMGvM0617xTMgDpxOHb2kUYx7pUppLKhqMYSr0CJ34DaP11zVnI9ykMbD
JnN9uKzwVjlMz5YjE2syzd/XhpGVCpfw3XSSLpSLDuFdmJAPNQrqmpUl3jFcSSbR
Bh6ZTu5/3449bUk2HVvjfUdf1qITi40tRBf7Fafz6t1I1gx4uapmJjLXQQQXZSVI
wNk6Pfl0a/ZNX+yXGeKI2MzHzvvMZnsafbKxIyrJvikMBzaNVkqyFJgcnUkDhJhb
Z3XHEZBfoEP4nVRzYO5yXZzIG2eLaDziTOqqz39hbkU4POolb0PRkZKywgEDnf7M
OMnJTLu1DIEsaMYM6NDbgkppr1ZCqU6OBliObhAA32tM1EyZAgKimwI8ZOx2HrwI
5ra30GDFDYyycGz0dpjLpsek/MlZTLWkCZ3mH3kfgpftSQCJIaSMDty/53WYzGry
XwF+lFxEkrUBq3+kdEJyBcwDfWj7yH+zbaYnuX3SV7u1Pd2VhhXu10cqj8lbrumY
Bo79lrLxgQnay6B9WlolfU8PTW+MhwN8Yy83Hlq+Tmc4OwySWNo6H2VMJIDXFrr8
AtpJea8QyeBA/j7g8OL+mYdMcfaY9HhKw8B48beE95Yr/l9Wa87Swq55qkdUVk2V
nxRhvLkkBAroliQWqLXxMRIPBACD91NI6O6Q0dvEZiUW7pTp99TC4aGfYsekihI3
nV7Hv0E5MIaspmQQj8FFLL8nWlvXnCpfv+ncoPr9IobZ2WzJqbrKXIiH+uEJrrR9
LeZu4lkjkuQ0lmRFyL2qfWrAgdFV1r1BZQn6sBQrh24E0hKQqvx9X77Q7SgG8rMS
fYwgN1yZ4o6A2qKRICPbY/c7CuR/09yzwtoC4+qX2JFRGRlsRhBuyP/LJAN3k797
IW3bYbrTJxMmCjrETRcuTNUeq2/dt60RHqVMTGB9q2GHmj+K01AxRU449sANazgS
8sx29Xjc8M05kRrynGunw5qpYXxKWIjqSuafYPa1dEw494iVS7IgInNDrbqoIz5M
KC1wVJp8cdYtL9TruSnsNfv16Vqtl7PTYqQHTFdununX2DkOwb2oibs53kxo8LOK
WoOvfyUUlOZlL8RbxAXmeDTqGIuYHZvcr0EbK0taMdDFvkCdRuWgZeWAaDa42mhp
U5NRQhAhVqtTN73js94fLQrc7h+Gwe9AgXG/ljxFa9BsG4S2cyovq6WxeIBLZCf1
jMIhTe7iGIuzCvHgIZBSrfBU/EMBevc+GK8M+fmZedQ+/uFJbEbNf0O1VW2bEN10
LoteyUglFhcR/U9Anum7QLLWzP/FfQpkxumLXuQLAA7qZ1Y2o2aCBawfVvMKjCaA
JMOYvfpboKQrdxc5qpW7x35VsAWF5rKTvcYrXx3UZpoguN65itow/Gmnh19PIhFZ
FQlGx8O2zOgA62H1nRfb8Wopy/tlungPVnIEoOhtvEmv6DdIQT+IwRD00OvytQTa
H5L+No1w2K20Vw/c7b88Q6NTWfrR3JwYiBk6K9v1SfbY+ajBKITVjUW2vhuRwzb/
74+/deyIFwfTh3yR78hF8YcXH7RBJ6lUc8kgT7xkj7HjSK1Bq39wluIEDJj6XEzN
A86gxgK7Y6EY6gn8gleCNEBmPkcfUB7FLRMfkvOSBiUT2o+ZfEsw+LorxfoFhk3I
irtA1GV+BFx6FRxrMbD32URsPObyOolZ0VoZ+SOHUPUxB3qRrt7VU7QWoS7BZsA8
MHTo1kXI4qROsxjwXRmKSZRtcXZP9Wg7sEgw74ozXWu6MWUkvGrYJKrJiAh15GW0
zLE2W61h+2lJZ3SQS/0ijbC1hCmKzRBOLfz61EIoNtrteKqUVbXU07S0gP0GvY7D
B9mevx+MUJMe4DBYM3irloYwDgyyEnRNdAry1hE12h0l3CXviW2yYt1eedH7ep4g
W9LPYOm8Bq/gPy+oD0AMCnIQZHMUEUiy+LbSrmhYvfwWb6kdw8zMNu/QmODutN04
j6eAl1HRGfGJuzDbAEe1kgsTSOrf4EGUJXLvIoe3sM7zsLhwxPrP+gP/BynKcpvr
8QSteJYf1HWMOV8K2tJt7ssSjlnjrDCN42KYfwmcl4LfKR6Vu2URfD916Oz1xyPm
ZIVU77lSPqdvY5sp1PwLBsAM83x9y26XjOA6USKKeJUQeF+57Jwt0DQQvTKGquxp
FZ91ytts0h3W/x0Jkmjo0OkXfKmq3NUnNLuu51YZ3MM1MFvHWeDs0koIMqyQrFDD
o1YwbU8cixisGOH069OK97jwMGTPCUIJyOaLO3vd/cX3cj2HUHXsY6dBwEezPOg5
gREFuSBe4QfED4+rzBVFRle0FAT6XDWmpnqvXH58STZCpE7YQapZ76R7l+5vN8rF
m6cQbPlPrYr81aw92xo3RyMUu5U8Qr3eg+5ZOJFBsv5W3TN6AjSE5MPISD/w8kSq
DBvY11pSSamyI047zyYEE9vCed2OIg6+fL/8CVgJ2YqcVU3t4WLC3gC1VyzWstQw
NGXUIkBK6+y8LDFscVSvl5BggOcL6NjHSg9+QxBslaYtYOggr5K8EyzZNrZlV0R5
++y/VTmpZBGOVxHIzwyk4KJKaTqcJ8C6ixfg5Bi/SPf8BkMwJx+cxmVCsvJKfTCW
JxQrB93k3ksLVzvJy4HDQ1TJK95e3jvQigznUSxM6egWfoNdwfvjt7bxIHGFlo82
AqGWkxH4wXySvHarX9XuU3SOPcZmumuX5V0lwK9/pf/wY/33DgHF0KEOc145x4jp
RiiVz+IAwYiWwRPdueC7qykaUEMvtLr5SAAuuYEwek/jOjgTJydAUDPZIW9/BmSl
yqKPrJJXoIqMgXjr3ekZS6nBnoePU1bvunKzqrFfMV4MFYr5Z6Lg3pmVOVD+8WRQ
SVTqL7rzP6/AOEHKolkVZbLEY8TalEZYrBf51HM2YW1/qyaqQWYIp06sMF7GzrXq
wFSGf9HXR5Rf9NqQOAb1EwXiGUNTAcF/h5ZEpyhCarFRVvMJTdIAzFga91IR4/cV
Xx5yQ5ckytfkKZeUIYbHjR8DMyW7PHBEwDtAxa5zbhRaQVT+K+OywhvJx7Z1R1He
XW6UoJugNRAmtFeUwk8oknxmPrlaJawaKWxsWtEsqFHwkD14sEQwXlldJ84ucJ7K
7seN5MqUamW7z2Mokhtu+z0yHtloJRaQCUf3Nqb4NeB+pYAl2z+f3zcbGrXww9KZ
2MIQH3tSP0nA0+pdvdybEiwqb+vBSydh2hka2EtW0kgz6eK1uMdhyBRubIhjRyPf
IJu4J3buicTveQ91lzOSFlu4JbHPy9ytY3+MafdQo5nHq2QfR77n8dEu6yKRyd66
onNh64RBwvnZq7TNTh7BBSM0bCTMNKLrZamO7T6HVdjyJFBp1vqNaaEW2cKAY/ml
Tm1v5+yGxSexpNygmcGmr4Q8z1aGg49SbAoV369azTAu8TD6WxeCz1yKOxRO/CsL
esRUScR+f+OB6kbDQwgOkTsd3Yi3dZhWeyNwY++aFHJLJD1qxgUsxVi7Y1antGUD
IbrwUslc/EZwO3IPkzQwy9sPGXbbGxJi61oCWNjlv8AYRdw0SqbwU287i1/xHr8b
BQc7uBkm9Gsg2+KcdTcadjmYHCazo7OLFy4e6dQw3yTj4veokiMCK2qtg06SzQho
o4Q4V36dx/5AhP1iIT371H9Q7Za1mV9386p+d22x0rIHmdgL2CXcb73zr2uSTgG3
bwUTAsXaPSvv37fOg7iYqXM7yTnuLV+qlbEPrxQw7PRNBcGrIyDnDITCHC0KiMcR
0jTgYMQOCEM9CMRi5nYs3nngdHN566rSrzLdRAFkz9tykacqqQ6PWXTkk9R0MBBb
VjDeAEc+ViEbjSFSnwp9U1yUYRAya8CpvfXhEx99+Kev1pZYAIepkKfjOojAmBKc
djhJlw1pVsmfhzGGgMEf9MdhIQttdwjxZQiqWhybVe+YYnwTiGQ9DFa3PYsYiDM4
ZKyeMJWP2NN9Sp38vDbuRVVl7Eoj8k6RzRE+dxfIN//zFMW2J7uha8xC53iDN8zx
yBgw+6NHXjW58qjhslG67GPD7SfZ28Qe0AKE83LcD5+USgGOX0/HQYVVTSDUOW2q
eAM4Qx26YzZFuaGnlpaX0Iw0oFCaBAoqRAPpZ5SsIwrEXtKLXIbMLp73iTM+cG+z
H2/ueb2nUib2s8l8NAZCnrcktA5vEbvUGjr0rCCsugHsrZRxQLe/+1otBJIcnf6P
oXXQNdB/lWR5cvDZ4Jk6rZSG+wm4uCasGb974IK9Sh3Mx/wSNuQ/RL0Ob77r3b1w
QDLi8ElggSc7Efn/s5J6C1It4XG/1XBpPn42yznUUdHulF7ZdVSig+C179Y1Hq7d
x2JRYEJoJXEe3tiDiT6u27i4kcfOC4ELpuVVFS1tWRYV8byfYx25OB68na5Cam6Z
szcC+DbdpPqmRta5VbnI70pSMH3VRfpHRWYUWsmbOt+qd4o6iygZ50AoUtYB9g1p
iXJA8z1HMooAI1vziUaIVQ==
`pragma protect end_protected
