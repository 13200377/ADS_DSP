-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
XWAvhhb1hPILQ8wW/EYsVtLdBevRXc8a301uyszElONqEyzizlUkF5UYOwxlUBe5RhGBSrAPxLbi
gTnvmX9i+LRvCon40Y/JgSeZmgsmORvwuDqvLkEz2ch84/NHa51FKfZltRCw3mt1wphhYb5wlL37
N9Zo5ipv0Qmb6vLpH/0swgimwcQAW//Lm8qLapOBVN+Aj8qN5hB/qZDKC9kfClDCD8ilFcwdxjoL
wGoW7MhtuzeAYWIpc2Q6tj67oiWoyi4L4sifORZmqPv2bCrOKCUPp16D0ghS4NMyQHQe2bqE/nm3
H/n42mNKaF/PfMONgk/JFJAJZSW6UlsRMpquSw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28736)
`protect data_block
ZYX78PCffPIvSSqTCh5Nt9NSY3K9WbMCdE6RoEqB7HAIR29Rc/kFe9Rd+Ouee4viuQGPk6HS4VdU
gDR3aeHuzo65ir1nCsGl8nMUyTihnr588QWGL4uiv1FJsKKMfXxIPXcVhXU1879dXY5QgmPuN9Fq
W6hljT82Ulj4y4s4wvdP4NnvFuvfGmYOJA4NbE/oieUkgEJNXMUu2LFSIteSo/ahhoxifyPjcj98
TxDQqduRfvR+5IvcNDUi+sM9vL/8E11v1q50LZ4Sx5sQIr+aAnA6Cn2slnKZa3wZH4Bur3jLzl1f
slkFIBFZDcDuJOOeH+plt0H9QDXna9w2OIMU0sEJglYsE+gY7T81zIu/kImAlyivWsx0EAxSKn34
QJX/cAKUU6XKNOiBFMO8OfB1bWrU80wM7G70s0Zyf4qEJyhlLkjAUWDUymg9B6cZ+aUjIvFnK2ns
hr9FAg+IikO/oZK2MeRXHU2EftPV6edvxvXcWvHavfGQtUjUDvyjC4ygFOcizxxTk9kMlWgV4sH3
utVnp61IrL/bfFICRPDNzRzJltLLpWoQGXr8BiaY1tEA4I7jBAn9s3tG6qEiVWrpJPJH/RfoZB6f
oTP8IrQozIA3mwi6jmqaF3xB1LkQiSU6dWcHrSeOKmPceNWXJpgVrqsM7ddd3slu+Rucx6/fSHc1
jfQIzr4HwE6PS7J15BafS4IZrRKw2M2XpMk6dPBKfZkhcNhP1Ek5o8vSM3javHxhtiT+wXDWv3EV
C2w8wecrNjGfsYLLhHFxPeDqWB0VGzZYXAb908aKSykjGqphM9OnxIfpq4p80ftOxleNs1yayhCx
7zCuZN3qtbo7Sy8bbPaIIUIPaDbhWmFStirLCARjxABe4Okopl8Ee+4q21ujbsE+1IYih8TN+8g6
sxsbbTO23RyuaW6CkzaKpAAKZfOvF2sT3y+ZnjohoEAmajtH3TpM8G14G4MQ03GZ7AsU2jGF+WLL
9SedAf8AjIAXqs9y2+FZ3O6RzUxCiy/wWo5AjziPO7It5HTZ/OMp8XumPQx8YxvBWfrrk0AV2dpJ
mVikMPfhYLuGUkPsLV2uB0x4mxNsw+l/XrQdOLCRkD9XLJzbjr3DKvwKCxeGVN0Df45hlBTG5u6Y
ZLpofn4Ah8ieDFRp/GLlqZbno5m22guE3rcoIOB2aBMwiG0kDwaU5EMpGhYbUg15d9P0esWLav3N
QUvbJGyPcmBJAAIkBFmd/z5OJTb3ahpTbcwyBP86K5oCPdOhN1ENVnIQoFh6T2GMABRVyBd/7I0j
vwq1X6gzo0SgRBGdXzMJLzmY16DuRW3ImQPLy4I9TrFhmVqx3mXOFJM0ivRS7dFTsmuREWSiTvO9
NTgaHvp7o3mNnr0l+w3NmfmeoxYGcGy/ShGSQZhbHQdykZo5+U3yicPN/prIaKonPQ7ksgxCUbj5
lO+pReU+zdKkVkv7w/fl9/0zJGRpd42iq8vZhld2xmviDtii2OAqDZl/KZtrsLSvzIqZYnvfmLRW
peK5tbKEJOxYujT9POc+vg02d9O49kRLuDe6274yBraKl0Mm8hg9YMNPo+JTEnj1po+yxpZrJTgz
VmvQyJRwQjT75I3BItitNWqoIRFe0Vb/hdSiYJTzlbbUM+uFjy9OSQpwXcs6xPYwNN++pf/u51S3
eqJa49Hk2zN4HEJhL907ezriO6Ml2mKBwHl0lZBNZg5VDyNVDYCqeL8stWFeevJKOfx4sROtDzX0
pUfrfCw8m+xckhwkpw5BvpFu50ZpGD7BukvTwqP10gqFkQ1SKaw+uK0Wx5a0DCg+lOMVGJKzDR6a
nLuI6RGzZzZ24J2U1Ohv1MBEHgAtoNAiMZRd30fSkMycTZN0QQg79VwG1AhJynIlKMAhi16aw6wn
6w22L7Jmf91jxw1cQbVerMsK8YqGD7je4zRpqm8JCVip20sX3D5xYKmCAAxmIKwypxeuzyoGI84/
XWEQG3yx0xK7z9+/djxsupXAP/l2VZMJboRpw27DnTlp3/cIfVgZ8nQl4J69Jqa+hbwV2io97tQL
DUWJJQZe6KEqBWBXis4RE+AUky9rkFiVLOzO11pBdGOZqnFj7ezrIh3M2py7vnpAlbJX3RrOK/nj
LTj/Lz/ELnYNwhvt1me2YD9ToszvHI7iklJAEvuFj3ssx2FFrBVFJLtMLJ6gngEokNb2WviKrucI
hzUF22pLzb9cVbgJEZC/y3SZfwIh8geTpO7kw18I5pzhrkszgJH5gtxx9pWHKksGBSKOeQwVZ8Z8
HjWiDlzlBbozxDcevMQKqIr8/5Fkg9i4YzPmgkDe++YFk10zHxMLPY76R1rE2FtZbdYSM6rncgEU
FdhBprbJlwXa3IfOZGxBu9rHM+emJt5+ewdFq7cliWU3O+ZgNeAJ/+6tLKJ+Gf3DjN3+VkLT25Sd
3Utgg4Tqc6XnKhkPwhwoUVEzaA2KV5Nkoo2hSSJaO+CddksiP20xMKZh3bL1tJ+2ZoY/sbR8REsc
rp1ifCmhTxIQ0nv3Hm/N91y2I1X7IzWchzx8uowzjgPBuOIw+cVfBABFTEBg/tFKa6Tbgvyo89GJ
MYgs6Z/ftULoTdtiTrB2psSxa3UrtzsQROTd4gFRmVej+KjKgtTM1Wu0F54hJofpGk6tspvkWp0p
CLc2k2cdcIF3oCkwvGOMjuVHNIwsqIOzz72YAOi4PYt2z9qUBW6ej7v2OqiyjFIzw9p+WUxZ0Dxx
s5u6VwKpX5kNq8rbKM5RyfWSVwH4z8ZM51vQShMbZ1P/emjXy89ECJsjJbv1VPXC0ACLi6eVQYUS
9PyBRBeYLNLFnlkF6Q455v5FaehuTobSaqAp7zAvQVyv9xjWNNA344lNBPK9y1qA/HUrcTwwDdum
JIXbVFxWCg0511Xy3nFvbQ0g+nAByP9wq7/E+cRJaM0fxBGB73ShOQSSZ7RJknXRwzdzIN9psKQx
A54F9sXuektDzQfHA7pOYgaczUxSUWdT2eSmV2kgpXedseUmttWEUeGNaT+VNC63ZT1E4lmX2Vlo
GL5U5nDA9hADrKAAPxuuKFeo6PwejNEv20oqLeCOEXh7WG02etTq0Vvpqnj79pAjsW6EWATH078I
Gd6hF1Qulgt/p+PRFCH+TMsXNDwPK74tPHuQcH4aj63j3Oa6TGFRNJMekPdKtTsCOi+hf2Jwr8vE
LZ0nhxjiwN7jvVMXp423CbSzAqBv38t9+RzHKYftK7H2wFfScC3vWUKAJ7K7kK3DDr/yhimTbouR
cLyvpKu7X6w3InFI158FrURkVcjBnmmXVNS/1EgRWqpS6E3S6wsjy1pGuWUwPYoi1ruWhw0b4tkt
4UYsB+vw0enkvG0waW7h5Tz/9rDBFBwqAFYuvTx4/noT9jlRbxWjJ06iYmEufavwSGvHo6ip7t9q
sFeGZmltgLUsMaedOhLVXZK5ZDrO1UKA0G5ct+9y37NDsL0SuYzUcQ26ZXxztvsa6D+dLkG8s086
YHJZ3rc1iSiFzYki8Rw+4yT5AHOOTNkGXD3WVV1vW64BokSYVyzOwaFGVvgqfrq4Iq3DJsg0sKRf
NIR6KQHm1D/5WK4UOlphTTVZfZnmM6EBXsRHNNzrmKgvf6mTDqvy7rX7bZGq292URVoEjnj0Cti7
2oluqBdHxDfeFV3WBwIMiJRk8dowXbILQBJxtsK8kCVWDE2xEc2EJt0VB07gq8tO2qCfqW3oqClx
asOiqOTPgs88ph4hG5DENvBWKZfdagVDzaT63KdsfLO2ZIosMDEGo+pyqkB6BYUQ2LHiZyjIOj3i
NEgqBHfg1mgCSxBQ1lRZzfqN/ffvqYf0VNWOj7/sSuhbB2+6wCZVVgMkaDzjmIiO7/IXkC1DbsrC
Gmr8M1nkH1Y6anN0x7x02wlat9FKWZl0wZ3fFlhUdZoB06DFh5O8md8fVf0+9pBGMI4x2+lziq8p
5zpyhIIZErM37k99b5MhkJc2yGuhiu74nFNdJIv/mfG8ufOqVaSzmvn/ekGXp/AOrP0MRJVbC9uv
WZY5pjRx120B7Qn1bqXGkS5fPX1xYUfshHkuXkpbZY9KIXboboPp2aWEehdlEWJj+wfszUhVNNLl
yoCBlOWP8ayJ/p879ZMXUkstu1S4lKk7aQcTKJMV6W3VGltmp08urja8owgTG7u1v1lkqGktjZP5
MGPO66w/oRcqjfIr7XYL6xqu3ddN3sQWbKAnKYHAd10FyNb3J1sNsdeIJ38ftKTePfmBpzpi0joM
cShxaTJAI2IQ9QiVVVoeK3ukZ2EtVyK0As/b1Hk+Sw29xYiswohBKZ+GbwFNIU89+3aOuD0YziWi
Ks2Dl37L7UO67aSwdtgwYRK/mCOGPEgE7dwZvOXO0fiievDcjAh9fuHyqQrz6wW6cRalEJ3v59O1
2pLesnu0wr58KCGnbeYxufjtQRsfDAivfjkmMLNELhlvjPRo7H38T+0s1ZkeJB2RYZ3kxOgAo0Sa
gkPue+Z3OFEC0GdAOoQ45evz/BgIuXAOdzq1enRHDSF1MEr7CanhBABlkphJl66e3cQrlDb1ea0v
BvXJML5w1BBBV/e/Ce6wVD6Zmk8AbZcD5+GYeoEWuhSLQdk/IHRivKk8MDQ4dewA2WHgFw0Ajucb
xNHj+K664VlzGECZmXpCbf+sw+7s/BXVUjaMqX38qM6OBxoX/X0DAJWpZZI8Jk39/DBB89DRdh4X
NursdEPRbABZ3K+4OatroqSWHEY8iY9yHA9zy/nFI5nh+rNWwS6Vuwj7EE1Wbx4HNBqLBGTXFr3R
R04ohN92VWpSbnPCG9dGj7s58OxBUBrFCErpD6FWDTwcZ3Mh12b6tD9xFdnW0egZTPBYPgq9bvpq
sMD4urWlqa9BSRDi+yxOQjPhhmYs0TAvAkvRtchzBAXvO+kNeLO5HTYC9OCU4xxoV3G6lXzlQGkz
0yT4mhpbV7zatoAlF4Anh5Cigb90W7b89zTVgItiGbjLMBJSENDnGBPgKZc7mlprRX31Ylr0TQp1
c8R2glEc3Y4CMbGhMhEFnR+yC4LOFmL5fHz0ek5u0Tzg/ocIl0nwGpgYH0Vyf3EO56F9ocbpYo8m
V1At+krmFSgaBXDVUkXbJKgx1PSWunLa/kxX0orrom7in7F3X8WzTzYeX+bk7NlnSVVt8EzB/ET7
Q6MmA4EiYdvGWOntiLTNydTbCnsAeGHbgy1Mp0oMh7T3x/Y6DHOn0wR6TgeVJ/l2QzreOLeyQC8J
raX5LRtE0LJq4jUmB1utJzIccaTeih10CTnabO5frBNl2xYKAKHNqQBzeBov4Zf06JbJd9yoPv8f
n1tog/UWX8moOKe7LJ+8iYbLzbnbnAEmzNHtASxumCqEHmjycfYFnyTk2Ou1/8Ozsaf1qcxulme+
WpM0z6Rn6xFD77Wz1ux8xG3ki8Kf2I6oVOFRYletakRMI0UG87QZbscghXeawwl8gUOcyCc2v0MO
jCDLObCBMPdRN8kPBHjYOSDOqCszXaHGp27Hpijg4nYEdwzKCactxJ4tPLnEshTTa8scgnsqGwn+
AZcay8yhXResIdc/5wC1w0eL0VITUHZFwMcZrDghtIuaM8Da2gQ1arlNV1wey1cb43DZYHw+mxNh
wTj3z9EY26IxxkG3ao9NydoHzZqvHg5VsV0/f3r9PRgL9GO0/aHfPkV3lVkRcj/zwrkUkjd07fWT
HrEyKZ6JWPvy2zmeDvRs2aNwdIOQS3fTxpRfTfFlh/rw+kRp2YbYBVrz6srIlWV114zC03DopBUY
IOiIZKH3K3XxD1tR0QNFkiSSO3LjySH6naCsonyCQlHWj+JDvKWlIz30+rBc7ZhfiFJkqlieYQKp
+TazyTkCM3y9ZGkcQ2z3zqe/ZObc1BRXPYNZ4d500zxfMgbPiFgfb+i68BfNAYXvPFFxvRdQcE9W
DIf/nNlEwqrKjaGU9wDNKiuIxTY221ZcuGAxRgdLaM/+DOc87LSDseQ6tzZi2RPCEB7f1/kfzolX
iKyVHyCaqXQL64pm5aCBFygHkh/d0U6YPsE7G/ZuBRAt1kI+DBO3K8G+d7INwjgotozVeoEDRDw0
8+BqmIYVbPqIUbr3hsbkrL54QPKIMrCfalaR1JVC/8nAIdKEld1rsjyvrFQ542sqlTeEhgcpeaFt
dyNXu5OKRy2k23vB0FC4SmoI0Cm0xZvAbFkXVOD9B6zF6PQIYmcPERMMnumjXqbEQYv9jLoFusip
Th0nuaA+UXEUERGsESiomYYYrAEne1qj0E7WdNq9qCVIeieoDbAsAfmkoFdd4oeevBHCz/eTVOBk
7QKO0EFrAymq3Z6SBwpMrXeTRdt2YWstGOXJ//IoYIusx+y5I1JT4l+3mC144haPfBd6iJEySkCp
rWtPs9GZkezvb3deGhrT90+qav3KLI+WI2A70cC5mo8ovQvQpT9lFKqdi74ve6yAV2ox8wjUNRQI
myWHIXa7rbPsa5K1hV8ELzhIPAHbTbwLlOIu83VWfEp44gZbCYQ8SzB9/NdgEkzCrVIJhY5TAmkC
Uwjxm3UNdA3Dm/7ZeFcjUB4YXZrbrWhuRtudtjQonR7LF3u5eEqNszdCNNsDxO6zbiO8fp6NGQG7
kOEKVBb/LY3XPC+Z1AK1X2sNjxSUsnudJynWim7vQSuLXszL+wqgHgiluj6/9utmAg/VmQQrZjkS
1FMKyk9Ew1OPXFtiznSSPjfQ6jvvEIqtB79OHmZXLGyMViQPcQKuur4xBIY3HQTXA5fHSRQuyEku
VsExXyWbyOLziUc307niOcJSmpT2yLvJzvvXa3DOjnRxJOmWLG+CJHggWVS2AXB8WLIPlNotjiW8
msRUr9et9xPwpufoNJ+MA1aq37yJXC8ulyZ2QSWoAErN3EuPuk9abUtvqa7FxTmgcxaQRhJGdmyr
5cnbAbYnmlfMd4SULxVWGicwqpfXjQ6YDiWAgZvmmaVZPBPy4F25Z3A5+0IKVDbi8LClv2yOBmxW
zomIISC4WbM5c5d/n0TMgPLSX3dXISUg2btDW04wJGEJtKLgNZC4hORSPZX347YBDDwigtNDdzgx
2WpFZByT74vjms7JG8/LxsDxayHEYgy3FTkuHQPk4yythRSOYen/djAa5qAZIjW5NacLDMBBitrf
7BS5+7xfOL9bSNnpLrz3767VpPORVJA1jt8VgsRUAPCqbe9cT//u3Npu/oIMUJMl7/krDYS071MD
Hvh5tGlD9hhXdIPMbEQ+z2bN7nknQJFdE1QkoSffsnkpTePtY70EXn9pEgobzqPwNVFjrLtMWJhD
T/UrX4ccQIAKFBI2nqtGgri6O9iJ8UI1spLIBG30aCmLGHVWptn++9seDAEPV7bIXMGXzYAccyQq
ux3Dq2NTHJ+/Jbo5gsv9YxGSImEinXQ6R2Vzguz+8r22USk2sUNBGVQvmEXp9sAio8ix2z2quk3Z
w6Q1ii+m8JKRpPxiqYZMHrQ81fosOpXzyaVzJ7ZMgGkYob6tr59/S9n/494fvEfZ8fzbEH11DTH2
oxyC1hQNGr2CyUHSyHYPg/5DPQwFVjSRCfqTWbOYU3e3TtHu/D7Fa0mjsLRRtmvkIWCUsnGZ9/ob
/vakk585mX4MmHqfB6a+iftpAqlziqI9qRmtnYneali2z4FMPx7aGDXMv1Om5pBGbIFLQEGDX43h
ASOs6S4S2Nx6yb758CnpU26WoV8AtWh3xHNGFHL1orifNNkjNmDFXcyJu2MnrEx1+3ZDiWS8qaXt
qrTe9M6Inw2Tpb6RZNAr/fD+N764Pgi3s5npaRq3uYgNW4D3RZl9WBvYF4aAp6SeMLZ/RCLdUrdD
dAGRQLlkvqFcivbgWmIm8C5gpiL0RstD61TZeth/YKCQMLz/FRKi5oSps1YM4fYS2NsT7HTpYFrB
7UAxCH8APJcvUO5pjtP4TxG9YCsMPO6PaQ9ucsZ2bHpZYnIzzZEQCGqpw7j8EGy6remDzBFmDRXF
Oj8I6LdLEzn4vUNKsn6oNbw0vuIUYW1xt2FOx5MsyltTpdq2p4JJ3LGNr8cZNpBSwFXRSO5V/t9j
4VEYKrvslBZt9iiouehYd5SulBHKTRp3ECZZkU4lAkX049LBzaVi6EgdeB62rira/KvPMyKjaF4Z
gn0eYk0lWBiVJzGgjhw08THmZc7jpD43seKmIy1hDL2stmP/lR+70pjRfAVvQMkOOAgxCzKE5TFV
zc6K4DpcaMTpyWZNrZ6NsB14OWwARFlO5z/vaRrXD0i0pQ9u6ZmSxtrsykIFYzeiqC6FVsn3wulr
3vGFaQQuXZ0Ejr/R3RhbUXJG/Q7VQnK+e2Z3wwic4mhk0rto1lurnYzt1ZAKxuEmE5HcHOKUz/ub
vTTY2QbFVtKD5jbto7v1efWyywxrmS9FtPpuaOdbCxFtZpsYSGe0Hbltm165sgCoUMB2KAZPO/Kl
1HTEzY88BhvRxRAPIAJbVDPfeIdFhni8+73BPWKmCxSwbWtVNBYCZ6JOJSNLfD/1RNFRqhNnTNzV
tX32dTu61CeJ0xGiHBD3A8Uz/10VuxobmtLMG1wF/iNrl0tteq4kfOajum6krYfHnbAsgiMA3/0o
fPSmnLApfakhIeWoctcPQ5NUjKOCWWCN0dH3wTzb0nRjEtgHV0h6KQnNv+JAeW+p/iYBoGe+TpbS
Oj71SP4cla0yRv7RTumnXHT7Hl51ox27pgz/PZIfZrZiKO1FvSyz+PwFwMthIFpraOWCK+wfqy/S
1DrnoOVlIFupHcT1n6SnTmFO8FS3QfHUZKDTQ8Eaccb3cc1YGT2ysMXw/iHrgpedD1GiIMaBWL4X
hzqoYhjNKR6pJ/7QN4NhPAomTRILWyQjimkzu4oMmepXVC6eMIwTIyysGMr8LVFyJwQhM/BFZVaV
Wf0IqBMLXnD4zWlLqZKk34U/7r1gl2Jj5EgBGCHVHbA+hCyWgcTi0mk56ZtVIHIyh94RBwbNl444
qYnbLP88REs1Dm1qdQwplcsHZEbiDVqKj7AUK21IfIUlq+i57rhO0F6Ju1QGpom16v4lp7ty1Ko+
fy6XF5tLAxqnad2LZxp9/g1L+6VsXT6Gnov/AaIORC4XXcUgooW2s7XrvNIRK821K0v1XQUFFywg
Qv84D2I4ZOjmK7zo4w8WIAlNjVXWQcc6H3TT2T/syMdZp0rzT/9zsYwwpoygh60VWrNFPXp+0zEp
J45upgMqzUz8NimmCRXG5TTfZ/v0V4YyBwce98tp22ho9ArVBHQJ6zi1d9j6r1Jh0OPeEBc1urnL
9BYs3ptglO+3Z/iBksuZg4zWBcpvUBgKlCj7q3SA0vgwCtPy7g+TJByJBTkSHaSTe5fp/1MiZnjJ
KVYceOogGfZPk/jIaUIdSnYRzO/LXdQKt9ukjsh+uAuqo6Fgr02MXqk0AmCYbTEW/pUDq7uph0mB
CI8sND3yZ55uqRry63VgZVhrmr4y87BVgvHiptBTE2mtUCKHuZmfHDesUkPhgdkIrB6JNqymuOqB
aH05WLKk2ouq2eAMl25UMOwfdQatg1J4FEVWz1KmYDGtIS8cWORfcZ6xLk9UBMQJTzkCwIZMmgan
0IrdpR//1+VtOSh8/wcIXYlyfDtCzgLhtb34qdETQhE5QcdNh2qtd69Hdm6N8yEiS6OarcCWaa70
ewinvr92lZgZT25aiOs5RugwxRTFWQKkcVgN4IRPPhwgwRfhvRfgz+jBF1gOz+wgKpZsyqOyn5Qr
iPhTPtgSE69jXIlvIrHE1LQlaHqiq+CoV2ZVTJTjI24MTGNIPXBuLX7Z/fac/jV4Lpn8UNFfaiSq
AqyfamDWO99R/WNQSgfzBdoYY7yzib6w1r6UqdZkwuFwbseyOIaZSaRHu0EZ2j27+XvpRdWP6w54
TGtM3gQYG9AqZmKqpkdAOhjwldMAhtekMQoBIYVyLbUgtpAMR+YyJ2nyNApxPTP0Vt0CZXIPVoAR
22Cjv+DH4ML9HGxG23AurwuVm5bY55AODZtx9Jd3xYiPbfzVDu3q6cdub/re/+s8dq2dU1HgPwV8
d08EQ1Z3NudplOr4mUZiZ70lx9lOQoFjdqohfUas8c/+lz6r6CgrFvnpN4lm1MseaemBFhlJbR7p
nbJI1kF9UiNDse8HxWlklHhmRPbT/Z2cviUipyOdfZn5Hly7yXXNP+Hu7Qzt+VsmW66rSX6v7uTT
XUcqHrxHCUU2qEZPQI9YMIUzj8CRa18wNRGzjZ5o66hwaMa06dVCqhk+wKEN6gMWBcrttx+NBfpB
1bUjzM6EiY5WuWj7IjFTlQQ288hA5qhzUUKcVOOolqAk/M4cKOEsVP3zEui6NyGBYmDyfQ//zz4/
n86cywvfZFTRdq5RKA2XGwHeE+tqVEd+prmKaRRJ5Ec6P7B321ofsnHBgLV6HaCKZlgvx1JZl+4v
9cEyPlrNH6mqrEPgwMGgv6vniGkjLrcaD/asFdBuSuoLxXaYp0ndRCyR0KktPmQp6O8ufx6j0Y4m
CZCYWoDOgoSMnUoM+zTtztLrOcNVYWgBHpnqa7Ul/458PTdqm5gzam55DRNH9rzKB0VoyUTdNzUf
Mun/gd3QI0mDJnTaPCw9hKQKLPJr42y2cO0j7ygrUw9V7CzMMOnL4Ieb6GEdVAQXBJeFcS3+exJQ
2zm5ejBgk8s0lMIPBt1dwvMHjAi1dL08MbZvke20kFPdYkeWftr5Ujg4jzKogu48KPWtqwqhpTtz
RnyKIrJXukyglsYTrI8n//i2+KsYc6v0Ceiixl8tHT2ayaGSetd2HMmHWrQ9hDV6pyNS1jqCDEWR
7aTS1fhE8xGKDDUXSJ95OBG9UIwtzkbrQzblZc8eSqJVoDJDTKqqA9gwbIld5G/nuE7jYn761wOW
3meb2DDs1soMMrR9rt7WRWpDqtG9cj8g3SlqdyYnLcSd6Enm0coyx5mmHt7EY1CPsy0vWuhMXXmh
QTuIlI+tyE5DP8s3U9d04XGVcjpefLMJDIk2KGGQRvvd0QokXOB0R7R5aWhaievE03huex4Vtd9C
VQf3d2zGErAYk9ZP09TBJt+WNRYtyxIcLvdN8bEBOh6FTk4/An27Pnmns/Uc50ilM/MBv5BRVxeL
KQfzrYwbknVGPbld1hTL7VMyw5M/SkdyeFQyxnesB0a2QcDzi05Y5u5GtyYT3D5kj/DCuO84y0c4
JDVPtvIfvpI6zZQk2dzPt7b1u+y8RKdFrbVyASS5ugR2Eb7Me1PeGmed0SMSEkVBHX4AXBguCijv
atZ3KkzjLV6L1TJitrIudzKdn2nNdUy902N3RQXFenias1WHGroir+7sMFjVt5ZVIUo+AKVKLCU8
azkLcGz6KIgc20/DJQufNxfZXzh2zcQ5IfDIIl2G0YGsURWNkfURNGVc0PVWA8OKEU2W0U86prt2
S9bZWi7W4Wp6Raw9zSBgFIUi8EPjLZQbTu58zdA/vroEzbvjoiiuEbC+vuqRRwdLQ+UcXvA1lYg3
Q3Wj6JYHZb4lSyrzG2fVoUydZgTib/WwfhULS/t4x7u0eJmEdFdLAl0dC2jyrQVvgmgmUkFBHpVC
PTM8Zgp69nqOR8VQzhZKu32AJM3ftNNGolGjf+/dYR6kgKsYmvML+l/U/1u4BmQ3ZvpYaxaDLaZj
6XGlSu76YYPpw2hkyvc42f/0zEI8IBAFMab2ufmhiVF7kNe8eiPMuAEbBzQSBVk4q3rwkLyixwtP
UTnuvhrFZLNfbf0PDvED8J+P1aBjXsKvorUB0O/6jgFso/VBr/dEkhLkHhCKTobo1MfryqJEAv6g
oUKyilBcLGQ42V1H2m0x1wZl8N8zxTHIhsQ1LhRI2LeRJ+PjuiyZBEFCMPQHD2hBg62tmRZilg78
0jpGkVCZSKv7PDnXqM7hrnLYWfalEogomgY1M8gRsh4E54zAm9fW1nT9ac5r3L5+ecfQ6+jEtXi5
s40h2MbBq3srjfodBhMev0/IQzc0d1tk7J69vtZzkJSFg0eh92jT8gHa+iCw08NI7UIn1Ku8ZQ/j
lLNFL4oOlFRg3sqCzIWVCP7kEWc26uOiZBpTEhH1wtvzvF7qW+cqmK1s8zeWggfb/I6S2y5UPX2E
Ff6IlrimfBgcv7PBNRPD4WbiMXpAN1sdkOg/0oEBrW3vMNsHD9S0P++ul7GO8Mb40IJvlG9lnOdx
SX8HdHiy/0QYvfnSIMbFFvO/iv4r4P5MZpDXQmKnSUewJmQpCYsKNeZAWG4MHy7Hx5krt5v+llu3
VQ3olQRy+9/bL4ZhPJP3oVDQ/du2+STnMbcZFx8x/YFymBha5J5PWv2WPi+sXd0I4AXu2Yle1PG1
XLX33GFKJt2iis8gNxAPygv9dl7/hQ1lAXPp5H6s4fPz5NAhVPoLIEA66ff6YPTEQwtPxg/zmOk2
WokFyjMJvPwhnQWMfqIOKl2tn0IIVtpw5d/vGdPMJnueqqsuJwfTngFUpPYcnln+c1rGoOvSkI8t
5SyEJlGG7QS6yI6T9ldq/FPp6emenMtJ3rt7fZUfY7aEA35RRw2vL8cgCw/sIvbq/qnfid/R5/TO
1oeIfmqvv1WACfv82FpbxxfbHzbyULjEu28CxbiY4zqoMqr2CKdQt1AfgMp8wZRIydjPFZfFqiJN
pWnsDTKUTwTzhnAdW3coknPEoWSG/F9vSGRw5MFjXQFJ4vIZjzsNNE6oWEG0Yryzahe95bSXN+6+
2iCSks2P0dKKMzAZqsyZA935qvjmxQMsIRRXPsE/COPDH4Ac03HhQ8l0CqnDqMp11U3YLLzbRlJ6
9w49BpII9z9JOD8jlhshQjoTtzuVgIzubVMP3s3ED+uv4y5iPK0g9c1C/z7N7yAEiruyaubtHwtk
fdSn3jKokcRAcntiYImci9EWgRUqC0inQnn6jQrzSvlZFGyFz6gAN3gHWCsTLwx3ZIBCvV0GJ/AU
HyDrrjJ16GhWhUj2o+x1ltaQrsU2HzcVu5QkPman4Q+FvQ8EXhufGhltOAsKkV8xb3e5PuLvDzY1
ndIY9QA7UcXIr0sBk2s4U0AP40sVdvOpSAiswnSCv7EPOml9kd5DOP77IRit/c9dBK7+g5cDsFG8
JLMXock3ehidA8MQ/3wKAPrDRmb6FHGV1J6rI0C+o5agQhY4xRIUQr5z5LcD59QNQm9n7NU6uB/I
XLhRbcHvDv2SkHbWzEz43f227ao2VTIzABWaBiAxdhEInjLOrIYLaSw90cLfDO42yt1b+S/rUfzE
79boU1pgHN1F3rshudsb4s08mhHqrYC/mzH97twW13XFwE99Zuh7zL7Zoh4dOySVaHlZ44drBnkv
7sBAn7BhxY1AJ7QUcohKBnk3EnchQO9m0Z2WrVX62uMIDRlNaDPWoo/zFVWv/f3PkHhYtR/yQltl
Yi5oRQf1l29nYLjeLWLDt1YM63L6hg19wze7ICbLtQOmDXUbKkkJCGhK79dfr7Zg/5WChiCpYaXd
qpm10LxuSMvtSlSOmxXOGX0TedHYTYSEs1165Oqavp7e7hwckOgKD0SZ/mkVsrHRW5fzIIrjOgnS
leGr56QE6jbKsFVp+gaiR4J/96EZYuAwRj9M6pTBQxjD2tAfm5Xk2BPACl+s0Wm0gCLLkM6FjW0r
dfXl1e8FEeDC+SOEnZLjOlQZdcNydtUGRchR+A9wa3+/g+0RYeIXZ7OJGnbCQ/z2DYmYgl4JlLfE
wT2Mti5VeD0RE00OEiASG3+iVkiNuH4c6eLJyClsNZBpF7Yehz+7m+Np2JPeghFnRvE0cE7F/b4s
YVa8HIqS+EmxX73Js6lkxY92BYiLNT6zmZUHN/0nu9+HljXQeOSj8y4APqTWswE0qQaJAa3f/zE4
3BBDM4jkn6eQRaeOeEzPo4cXWVMIalhlB7VLcHzwOdTuH1l3eKu/+FzEvhvUvDqZmzvo1g3KPGsV
2bOXqVc6U7StdLETLFOw2kqeLXvVkpttETy8HC76oLp/cBmjVQwl01W1ed7kZREF9P7xfk+6zsrS
lVsPb++y4amrxvZglRGQeq39NETxfshiCUVoenzjpEK4eQ5SgSWiSbhe7oAYrWbSeTEVvgTBiAvv
SJdUtaJP9G3Ws9EROczONxeeSj7cHCU49Hw3CMmOHFDHLSHEIfHz4DMY3qa/sxXjFOeOFiJYZfI3
H7cXQk+eN9w9CKO9N1blhZf1GQUH2i4T79zpCuz0384BVN+MlqncQZqOcu+tq3iwL9UatxAQUM+t
vCLTuQ9kEx/AB1SJchvVlS0wJVFYBURXnc8Xo6zDt+WFYJ3UGEo/ab2kErFEkm7E7PrWHbMDkfaL
0etCmk5z3jiaIhwMeS+oN/I96ulqyAb9mZdQu59TopnglWGmSPjwk210+6ODErXpMOZMsVUYwRTn
uOQdKh/2TtzIXecRPky2d4Byv6Gbdjtgo+YUlCNRfJg9wKL73kIW0FOqWU+cBUxJkf+yVh72ovGy
t4ssxGaL5/eDv6EHfSDS9pM4JzHasOqJKl/k+2lWu4mFix/I7hHxK/iQd880D5Zi0lPq7Hee6VVi
c62D6Oslt98Dprtmw6fCiCGFTRgFxGGIYE6llJ9gQ49DYgIuMz0wcNns6P9gKRegY5trOEiV74+7
uS6pjEYB4OgtiE1HbnoFVz5v7iVvkFzU3LIlCFdhaEhXUxZAL9D2GM8C/2UWG0WbFq53KTHqU5sZ
tpdpOU0WFxS8Sc6pC4+6hOqAHGHb2FJL3Nrc07f4Vr1162QhJ0z1p7mqWiy8KM+VKb3MvifTspV2
6dj09oK2hRuTdzePgB9dAxXWfmZJv2ooGZkomI95zwMU3rkixvvbS8z20RlErvZBxqWbigjyCuzw
ccZQTl/GWcxnm6kNW0nEs32/wA91zP8sJO4FEJWOUlkd9mYhBckXy/nZYVfINpcaB0bolT+35jJD
PR7Rab564Nctz+hebtZM3mYwCyo3WSyY1jCa6k0ZpqFczhaXwKQZd0jfNcWkS9dDyc59IwyTtnrN
04qFVTJjE0A9gWGvYzmUbnf+enBSfelAxCVqpWyoMrwXjELwxRUoCSwPvz84x0X7SqZB+Ks6VzBm
KlX4trLC8STRjb/UG0qyL1KdBVgv7CRbSl1wG90X+tWZK3hLoFSII5RSfst4rjKYjjWc5EBXfJOM
g9FDgQfEl6JpqcRjLjW6OK8JrJaNSnM3t1vdypnF0EWbOVm9xVvKYndERqYGb7xbI+/vDpE/x+tL
afPdHPqz2zGFSxvkaCFRl9RI8UA6miPjwvCjHIedGoYBcWkYFbhjtbzKqgEl2uYl49gMDru1GVgg
K+jOwMv78nG+KG4XDkIZQNeZ/HInqr5Z+uKO3paYC38ShtlJmMXP/v9HvF/u3GRQgPg80eSG16c1
x1/nz1vUxgi5WghYBmefU6FhIky8s+iayAocsUqWaHZvfmSOgTvuCXxjOvYaEs1S+KwdwLxJpKRr
NIlIe/jeXydzdBtF+dx9NAj/wmXvmWOVhCRnZbyGVh4MzAW08M6KlE5Vk23OFRdOtu4hEbYhVYuu
jQfGWtaSzwkMQDMoSizQAuPuxy0LmguxaGk2DFMiS597QBnU62eB2JniShPw6Kj9lLqP56IX1Lpx
zWuwJVB2VbBQiVupYZXXcFgHw2FadvoZJqbAqL6Zg02kOwC1VYu2y7gtMlmWyGJBbKmQzSg5k8CZ
CtOrSf7N5Hwy7IYUhsRB2Rx2rT+vKZa+ukdhDOMpHR6tSLYE70rQnA6q2NVZGwv8ccESZdP6dToB
jxSw851PhezPn3jQa7vyt83mOc7HAuKtr4qmki/py/YzQoQfVokHI+t3I8paBq0AuokZyceLJxlB
N5IgVAOOq/QnG8BSznuKkfDQHplHu0QmXbnTEVQTSnLj9dZyeQ7PBrR51pw9kp9eosbmKHoQu1y4
zmrMx3i/JNteLZTlUkckDA8R7UJ8KEVqYeaKeBBvnKbrSnWSrORoXqFk9auj7R1Nz/ExqGzYsuUW
SzMg/HFIdV+CL23O2pt6xBSjnrcWxoMCRoJetKzHrk1vfNo8f0Bq0J8bMZMe5tD0CvXomnF7okc3
elvhCRrfn/4PUN5TaOLkr+pZkEpl3DAAkBZDYs64MO643WT4SA0cQgZrqf0w5vbTInFFiUYXt/t+
IL1UVW6OzFt0rTRKGnKGZ6wbGl+WNNx3jnyWQdWpdSow2YJxZ51cPI8x+i2fgfRMQNl508yNW+hu
Am8nCtfgrx2J+tH3NRlJ4tAV13bxGhM1H83sbOvArIc0q4ngPAzyejyYx4qjd9ScqG3LR+bS8hlI
pJ3VMPNVdp0sdOstGx9tFKp8WQx+FUAllM8ldDMEnfd3yBR8f/DShSiz55QTT7Q14bPoam+VXocd
EWqU7sXv4tDTU4tE5eaqdkLK/FuwHm1sG+BdC2kVKr3ZNgrVeoEsgF+VtxGI7UVEDW9heTQtPLKr
8AV6rfqpwGmiHCgNYNq9GM8tvfyqdLvlQyOzRf9xMfp2qR4CBfb0WKANrKHrizrxRt3ibi8MY68j
nosWLb9bBpZVC3CNEwt1wIHVS2xgQopqgh6ON/IS3dCkELuPLO/qlAPefyt1zyRZ19EwDEZ0sKLx
z/WC/VD7L7aNEW70NaVMUeg5Pgdb1yPqS021yLwMd+YTJZxcDpm7MwULS4Q1bLzM8hjoTCEVp9yx
9Sgh/99G/wqWZ9v/tTg3UWR8yqtsL+9yMUJRHsr5lTtTjrDhXIXGRn1/2qpMfKl7edtpqBRrlUwG
x96Kvcx2YzbpjrOa7vScfoJ2skY1EXHwNC72KBBMIn865gtQuf5ZsRi/DgrTx1MLg8eG4QCiUnYW
BrfXIwGRmX2RpQCnUx5g8cBoprpG7E7e6pO3QUBZuSP4W9TWt9Gw3lQIjBiuRU/bQv3QXaDsneP3
NIDXVdqhpuwq2pYbqgzAJuJyFSoL+XqdxuqZF83CGuCdCTfZ+7ROku8D7RMm2Px/VPNY0HEbxgad
RTxdFj+khxEs/SNjWugQG09kmMelKvwDChqVSTpMGK+ijQM+uNO3aeZ1GON3sEEj0zy+d+9+IdAq
3t7rBHQSsZQSuC4Dz4Y5RpXn5yav50yK6Uq5VDTwfMsImubHCTfuSxjvXQkPiQ9oZQpd7kZfxUdl
5UQQd1+nsf8azUoeSm+grcrTevYYqVrBw8BaVIgeuMAWW05qXW3ZiiPOmnMByulZ2IaYaTV0nNxw
7jfKD+3Ra5ylTgKc68gL+EQiBfGQd8Ynz05GoYUsmW3IGPQiKleBrkcOdKaKfV1r9CrdrXkWYlqP
sdtIJCEp3PEfsZbNkyu+8+EE+VUyDL9LV5fuKUCnRjxHtLxR2ngtkKZjSMtk9iZTaNhDj6Oz64cs
hxdNG8vH/ETLcRVSMULj6Q8eC3LyRDVcc43bj8oS6JHbvMfA6iZRH3EkXMwWpQKrMVpe00CGrkzx
gbsYaGbwystKZMlybUUU3MWezG5oMK2KnloWDvoosaCyd7YVrCdrzNHJwoWO4Kmp2B90tN4Q4O9i
/wLVtT/+/ITeZCJQpUnmqWYCkCeH/e3vvGi16BEoWUdS/L2J6OcJfn0tFjozWkjzRZ0jGTVNHbBg
/z5LtS9Euk8ajMbnHzuKB1Qc0Qz0e7NGLXYTYsD6VXoeEmKKhFbZren4xgDVZ2gU6MnWdxIhf/00
EQK06TChmR397rTPfPhyqf/eJnwTDbV6Agvr2DguZj9D3mZjHD3hMxZG4i65gF+kwZ9ZflOWC8kJ
UykdokfORgMfQfEA1f26vcEzUSRRLpTzuwtAEvnTeau9rAH1/90HwJWX1ZtGVh3NkedMwrqCQ5sg
vlh3/gCaM4ZK9t0ejLFqEbwCZmx8/oZ9pyu85TS1gdLZGQKU9W0gVU9sXrcPnccNAEPOSS9nn3eU
VNsasM6ur6ohm99KpiCMAb8H90eKhkCcwcLijG+MzC8Hr12dZjuiuJ4unl2bbQLHdUN1NHT4t30H
71tnSSF1wUaAAlEXW5Abt+EnmF3wcVSeRP4YfdXW8dqlqnFej8tb+MyUmp+NcCf384WUXGV6MoXX
AC+zg7jxCKRKHIvfD1Ygw6Bq0k/H6IbXf4G08MR9mFxYZ+0NiYsyR+aw3L1G0WScpgfzDvknIaAP
LqWC9IBsewbfXidS/dWWy9o1exdxpU2N2PmyTTqGAVkenQJBCQh1xF/0C55UfWohXjFEmeBAg6Yy
u38Xaa2Qiec3ec7de/H/dFI1CzW4WuzQlXFl/OfZyJKo5EE+Z36plW5Sq3R4dbGZ1q6bucSBe4Uq
XisiWjOpFnFM0aSCyfn54+avL76T7o2TWxIK/UHtfHtaeRsfSL+smiicbl0iz/Oc/tIfv9fFdEQI
jKgNrVJ4UC7R8SIP/YnbY3yFR/Y9oRGh9NQzA3aRfWd+F1RL2IptKCkumunVXykNhr4Zx2QCiNUG
Rj+3yXHB45tW4txLD2W/SCulE1/zmE0pOum2c4TK3xyWA1GUCBeoOIt7e2d/JkRv69H/zpj5Ec37
ZVYYNXvj1qbTLFLDnsxpwuC+tTOw43FWEXHQNGGfmiM0iHhvtBGXf5OQu2F9aiHqWz/rcmnGdW6W
m0ZnWvymmwJHU5fBYw0pk0sRcHwBROHPxUGoGgfu+HSkfqc1bwnD8ns0TlWk3mAP7NSYnOIiwA1M
mFgdaEZ1zxyyUNwH2k1PXpcwxFPQIyX1wKwNGJtpbBi1Ap9TvO4MnpoDhUfH0uo7C2zHF6A6hUvQ
hz2h8ig1Nj+j5VmuNsm3LVKXnYQ9BMX7BkZ3P2RBKZ3i7FqlpzBUK06hyXPWfR4Tp2TVltkj3voP
AqG8TaMUtZp6lkdxaDUGBvzw6y7g6pKEPtpxXNCXZRgIjWE6ZvsLUz3as2MJeLhzgLJYSNuLUhmY
m5g6F3/YvK/2FIzyRITW1RmPgSifATyfCFlxzBoCqlkOUiHoOzlOzMtPEo7fuoFF/XpldKmh+Xns
5hIJCYOhnR54wmYh1D7qaA+YPM5eQmv/DpuoJ5uAiMRx2Hfa72TMJvIIWXPKpvk5iPobD3VV4Ryp
UZVqFoJOA4n56IlRIjI6YPx1Bdy10EPOxUNTHX3hacO5OFWTo3jv7vCRSv+xbdUggeup2A2cHAl4
7hVdZ8U0gSTaSRRPbLj3nl4iyb42lMLsdDzOYlmo2ylfog8zXAl1p6v7IahIj7UVOsh/Tx8lYaUw
Llk7bAiq2oKAcbRgxAJ5NVnfnT+QQ+80IFG87BOg5kFGFRKLwpVf3h5bBsLeZOsOh0jXvA5Xcg/6
6ud/XYkFFv3AOi4lgqWwj7xwmupXhIcvemZa+xnubbplR0GQZLaAP9gxl7uvfhEzQnFXrxfKUFN0
9M30+Fs+4AF4MSkeF0mxbdLVJDPjMxNXOZxSOESxqCXGbVwb9gYcM3JCA6PJ648wsncHyDxTUf3E
AGmShtObRC+aA7Qro5zZy9T/14qTLqmAiuWDos/sKxs7MQG/rJ8xFsw1C12ToxDlYvhGZYQjnD2J
/OYapOutlO4OkkV59a7VbJUSWWxKMFJr0ftycYd4zNEKjPjkCbYFlRVRHeluCqis6UjNNdCRXGr8
koDgog8em/uRIkpCrZImIXokaYCZqwXgIqH8UkJ0gD8fzoxKwHZESFMxQf03yfVqgzzrtkj1aqyL
fym5oh6FEUC6yxjnYe0Ko4l92Ze6u8kF/dtl7j/dr1sED7/H0ME60cncNixW9ZN2r/zkC/UlYYJj
amsa6yVpsbDTCHMSDpPUrsMUk0QG33sFUbFGtVPdz/0ceKmQ32Le9nwEMiX9LG3UIafcDtjAuYS7
iY1WnPYtjCHab6GajAa3rfHablw2w1xKLEbUtPThJ592ovIHsNnJSGZKq9gXOfX1I3f1cs//g93J
aRVkg2vfr6mmKiqkH5NZoRv8E3hyqLzEhgpVKnilhv17TF8HS3RNMj3GWFOMrM3ClSqR8zfyW4S1
73guGYyraHZGk7WjdiEJTk3jFX3nzpDrq+gmWVA+pKzh0oK+kr+e2/SC2PXZUG33LFstjZ24al9V
kWTjt5Vcmfehh0Gst+9KltPiCe219RsSMLLXJ9Edd19FtQa4JGdX5zA+lc0OkIcjJRQYlFwuWyaW
q2S+27hnOcUNvgt4M/XRhFmgZJj/PdzL8j1tw4uVhudXMjLNS/HHD78r8bq4x7T/6QfKep/1Mr8t
z997t01eHuihCRPXdVbgvFYLnld29EgXuHytRoImic+wBjnqixsKxtN+pFowDnrkv3gyZkFoaElr
adpKbqZBVfTrlU/YrWuCvkfdjzzJk4hL2gREFbMaKjZ33fftRqe7TdQ+KVp6TwiZsPcDC2cgWC8y
uhqeNl8pStbqN/NlzOe8bw85cgi7KS3B/q1VTOGM9EQhtFapyvluIZAejd39p7dBulVfjRN6sKl5
N1oKv0dqoMPjLfjG1qsmLio6WiUpZx7WPC4IvW7ZDby/MRJsuLb8VR2aaKNjZ/3g1ovzUcEDY/fQ
z/CvGOjmFlCXKe9OLDH6SBXxkeuki7++myqJVbuQS9rMTrk28+ZRGZ4t1XLp1+sCP+N4De8ljZ4n
uXBfJ8VW1nn/GwnuiPMXneic+YcNSk7pRdbLXwKGz012fp1tPvi+rEIs/PHQiXjDJKVGSyG6DVy2
Vo12LqFT4m/YAmOVbQsDXvksFT/9ZWW7XjQo9oIGt3Y66Td0om2+sV4lVVq8JYr/cxPA/UMYdz4M
GlKaqd7WHg+0xmy3KCizJwn3zovtYWb8I7/SoKKxk78Me7ukVr4MNR8vxRRDXNQjyychRd5VIR8T
zMby3A/gLsT/qko5I3b3APPycNVB8Ne3Mbbrfr3I25M1dSAkqWTSvm+urGpQY1c85oI8DCw5aKqZ
60v4/9s9PCmBORLIhgIVykAsJ121cWhp4KMIqaSxDZOAOadqnW55pZwMXaZPDnCsdnUPX2WdvO7O
5O5zBmVKtO05B/g8JifqquP2+qcWLFPpi62f9j1rOUKBK6osPOphriG/x0jPVGDOmBzc5OBEILBT
DPh2uOIAX3IT2HF81uYCwriecNPFtrhwOcw3CrsYG3Mjr7rUh6vTMXf+iE0/VS5T/bCK7FVq4V5G
8mzdHNCfxSmbjeFj5qkiEgyUedhyJuRHOvW7m8g7l+LWgdCz1Svs8dE1kKQChy+7tJXZKHe+kn5u
5GNWxJOVUmiRH0D6oB9Wd4CFWvvVKEP9EoqLoVswDZjoDaG4fiJpinw2+jdBzh7ABA8DtMzmyMNv
Wel3EDaP4qFVRqoCXzFWUW7pyIrKNmNlIN8QzqMqBRz0bFgdHb6Mfbtkb5h14b6piqvRj10cJjqW
IV2Dp/3klO+8v52xUslXNFilCOagvmM8UdT90gWgj4A4WHlkNq6PUjmhJvaCoKre090yqfpMOMxW
BoraRBfZfUSS5ZAKsniwb64GZtcpk0qb+KT09r8QeDyrnJtWQUERQlR3epO0w0wIPw8lXH+4emsf
mmNZiSs6ZIq2Bt2fiPpLtCj30XYnanq0lCttube0rBKQRVTWAEvLzu+6K7dJACUdgloOFH/IYxw9
f+fhhbBpkR/Ki8embWjw9Nz6oPldz1x//pCYfYrxOCqXBAGAJGX2k+ZwUDj+iEQX6BLsuklhBSpS
gkKSlL9ctAugGwe7xU2rbBnhDvfEHY3q2HuD+ow9QmdcIaMv4dBTklDvOX7wA9ZcSMMSQt/VhopK
JqlqltTm7eUKSE/fQ7o9PRHO2zqmWvo0jWilkLE6qpFy7TxvWjrWZ8898ouNDt4ZxswsGn/HRypF
P1B7PQzyAo2zxauuAYgYrTJ/8fCWaPE6MASHs1KsGMzZWKMBnq2+StkuZbKDuPp2Vq4G4EhdzbTt
8qEsCDmVOPuXiFw5lWHSg6dotAkjVX0aohn7BjjSdK3A+mgQDl36jYMRUsCGNLWudgc23nHDaySj
fnD4bZcxKTx9e9EY8n7wrpxPqzJhqe3cyIDLFcSiC+t3i0QDqhi62kzlcqa8+5ARJvbXw895GMOM
e7afcmebwFzyYhtU+nAIbv1iSbWX8O0t5eFOJklpdzZiyKsWpzRhvLPH9wY4EkeTMB6eX66hdXcB
qhjcw4P1SfrtlW1Qw5kmt4Mz1iLMMLbXe+dGtjVVoO2OHVuj+ZctUcCUgZP1FA2IMbR9L1m+KY+m
8DU8NZHT9I00NhDyQsPwuxeb0HVLc1RGbcZcXXF4SCn49XHtgB+dpjhx+gW2nT6D0nZV/v6UW69Z
r9924VkdUqxrckD2pfgIKSSU/E50KSaf6TH+L+gaWm3GRwX7/Inr3lTbKCC9vBKCPMBoR/asielg
Jqm10s3Pv/+sUt3o1IkShX8+9814liWlgfK5cBphaYnxQXSU0U38y+McfwoRIyahrGJzkqdMze3G
E2qNJGM8IQz6V0ROgT4Lmrom8xTzNeJABWj3Jff0ndZxvqDM8nXAlXE7OQUw38caaalwhg1b45ih
uw2+QpltlWdrXvfigA156KqBnkM6Nje2uwn3So+7Hk0pQmvVWwaKOsf3SvpMwX79CqAMFMaZ/wy5
28rn+Vge1rjyrJSkB2htyxyDI473z2A33q8HExQD/hjW80tqfFSGjrbNB0M47alCDPkN3BHqJhdv
KNLk3zHIO6FtMquCmfOZEabAFU9lQFigKrHiA8CdTXFSiR7o5Be/P2mealiqo2Q1wzrrzsHsGdP/
roI5+4JlEhEafJ8P2gQgt5dqTNCMeJB+6eB39UudtqMrS6YLOvaHzQhfyWYJPvttR2BbLwtogOmk
RbxmHOpBp3IeisIuSW7MyQ6QV41sqhXbVYcb3VQM9K4poGnMznT4BY3nXdii4SCuLgG+H5ivtM3Y
CijdBDqaroQ0Pd3orqgPw19rL/k9hGcDxfy0HJPmW6yip1G5BeA4fNzpjqHdWH7Tk8LxvlrO6QW/
Sq3PyWzi5SN8Oy/z6yDCAbSkgQxnGjheDXuhcBIw2gMGnYbkA0n2+1jQfufMcs12duK1lanQiObL
qKYAK+5rA4HxUpxzHL8MVRAN7Hv4dtAaefKNAqdderF9vl9iB2f0wMhgJMWgluuRBRu1nWmTxzPO
qEkpwgyKdVgtZjGGZigxG5oefc3Py2zj5Tm2fPVx8O/o2fbuVMmyzHWTu6du7QCNQsDgRy70CDP0
UCfbhwBgPof8z/CJV3lGRuO0VtfOQz6aLxC2+Jg3rXP1Jd55/X3M7eD7u0n7BtqHEoXSfKwDQwCT
fOSzCe17bnOgUCEaazUpdOvZlr9EXh/NHI07Z6qn9aAByKGoaXxuJLQf8VqPxapFi1R2UzO4cGEw
vrOBZt8ZXiAcN+DE3Dwv2TH1zLNM9MUY0OVvROcjC6HjW6Ac0Vuz1O1qo6Vk1zQMPp5lc3+ydB8b
Pfuk9AoJSTaHV1yluHPbmrGhFVkIAGukuBZq/nvDoaWEewPcHNZuVGsXotNVDc4efUySlI6blqPx
bqUglapeZLMcMzdYFMtnuJajBRqz9ZsxJFi0cLJRVsqu7tS9Y0VBJLKx+3kGKz/bVq+0OFM+K502
zQtViBlcUnQIF36hRj1JBxJyS5xEvnTNG6ixRJ+kz1uPG/ssZpuszpYmECgDoR75limHWoMjZ0m/
StS4ph1QvtYOReIgzJMZghPkp9xetoeLNJk40irbRhJYvvmzn4ocHqBkarTaBavX6YQwp3R0Dyb9
c5qVr8+6yRNDdBYeCMrk6T4UqM+FUjZC+wl5IiTOMF+OXoCShdT0IHohgvWOwqiXGYn/AZ+P3gXN
+zR1sNKMJAtLyIlXrtsXfpLCSUPPrg18AW5U4mqBaEtqWE2eyMTRvzcY6TkUgddTPr0N0KMjv2fE
9vLUFPNmltsGLQ4IuPsrtmhS91InCx12365QpAIdZ8lHeN2ZekiKjQtfHa0aaOBBKEho84790yNk
wYTMRWSwZKB/piSbnIt5NTB7OnqPma6DfKPgvpqAKkfUTiyA+CzViyfPB5DeI17MGUaAv+TufpiD
BfHjWiQpLIzjc4KUQZe0+Er6RduhxDAbx/SfdhWjN2HKGQ/n56caB/D05Q5DncXwhOAvSk4G6eWb
noLViYfqbsuwFdocOPCJWVKh7MVLcGR6o7TzUKi1dyz04pcWxdamwru8C76prFqc+HxR36TEDJBV
fLm/0+Dr5mvG4qHoq5gJ4UuQ068+EO5RPmongmT3xHA0E2qkjmgbCJSBHo6GVXxv+CeqO6S++RzB
BsaxMi0vzvqpmSN6E4bKbqtXZ5yBgazvDWzGJY6sFE0+0RjQyHpgOxLq/bztI5Q3yUb4YtLampkI
nzXaSQkFsfuTNjEO3/Ze3/eDVQwAs0JuV4dsgbW3xiZS5Vcr1Gek4kRS4qQd6ApbaYSzCaArkwqc
yt1d1+w27OK/L1ERZBXzAb619eCB3pVrMLyl1mYlo8sMylk3z1+EV3zzDfHJtc6/ERNwBT+dmWy4
M79rr3Q9eeeng5CjcZw2nMzT146g33wetOQSW72fgfbQRqAeo9n61Qev2gn2IDfEdyHBr5CUmaIg
jlaTUHlOyFvXP/N9P4494s9dKZZBSzpD4OvKNjAYppK3pQPUjN4mjckZknJCKyoKsZdWy+P0kqBh
FFkCGHwPrkrZCLnQdsqEyOHONPgGSBOL62vaxMyLb/LnZlRmipGtmuXT9IpiKZ1WLY3ki6C32/sZ
JGL5GMrqo7+WmIzXorzuoxYPwP/PtsicfL+ARyewR0kK2hjDTEJ534tV077WYQ/BS9e7DswoNPJW
z3L/LyylUiCrOmSQxWQRm6Sfe4JTIfj0+RNNtauSV0+TFfXIkbJleffSND6wIe+bxgg3mmuyFHOb
2pHQemeqkC10frGcSbNKIaeesPhgZVnQlPPxCx0r9YesVEwnqi/4IJGQ2Ge7mg6/X2oYxwIrWow5
DGj9Me1a+d6VSTcVYmddL8huq8SuYu51el728LOmhzoqoTxbz4VKGDL6a9zNrgGAXBvvaLDyNyos
KJpGPbD4BjhmeA0AHI4sV8wgw0Gt9geB8fl0lKRuHM3lhXQvuNtbH52n1vvaow6v6uvZ3Dlj2IlI
16+G+hnJhnPfuUB1k3qqV/7KMldOU/iJFPHTZA2a6GtHXV/P0WjU0zqt89hEekeI3M2XYZuBhP+2
ry1dpeXiRYvHiqBcuBgYKRPgKv9Ok+1XYueUBt5+2NjAWsmJJAWqU6G9MXjxq63qQPRGPL7Q7RaO
aR9FuwzHW5SqMSZskfbsiOeyy4MZZAmBsPhOpRlsTEFcRhWotzAG7mwFkhaIWh4ZkZ20KG7qWYmf
AdViUp3u3VaB8j65RfGbXawJikrE5Gi4vL3K3tLWdnNH3c23iYu8gRlvzNaT8kh6O6xdSJFhDsy2
u5W/IPTisN7CMgtDVfqUhnFaztFFHb6ODA9dXfNNvFepk6syywxdh0/i+apmOCrc/LGpt1NoK/Q/
90kfEwXOmQSMkYLXjrTPKQz6A7uhE+vG746Sz07+dfdDrISv+lULC9KbbazwelTW96dlk432BAti
YNZ90JkQ9pTJhKk86DSo5pONSkyIGxrZBGfZG5x2P6LxEuCdG6uLzCKKVVQfZGQGRwJ88y/ud9ZN
LNO0nIiJkQX+HG/LxpOCAaf3P6BbYpczhHVaMDVfSvIxphSG8spCBS8tAZNX0iPULpgIBLrMa8yP
1twLij01NPw9oU3CpqjpRjfnwsL/+q5ai7FgHU0sNuwL9TSr8A3DAeeEI+/THnhpLemuh2PSUYTm
gwDw7rwW7APkurmub1Ntpi02CGHiq93CM7gebZJ66y1/aztqsEDAsKMe6qDdOalybP4jh8u8u/pe
4TGGh5v6drRqaQW3rwn3AnEhLimHVBHhLM2uSwPTJWrBBaRKZQerKE5zeIV0maT8ROl/zc+CYxb6
KuSlNrbktFNQXZCXZ7iHGDddptz/MTJgmQ+X/J5bHFDZnrkLX2cgTjUG9NBA72Yu5AofV5cqsMTQ
Vn00RdojHTxoIJIEuarAE0+YcCQX4pFymxEU8vwEqDnmdmk5KMvR4MrHGog6AE0+eYD2yiQJYNx7
FBuSSVILVwq5Zby2Ecl1RpjE1U4qMH5R6GRyT78oYt+EmjNY/zg9E9uoLLclHOHnPlyviTE3Vlkw
UwSsEM10QMoP2CZkb7XBhgwX4YK3BXVf3mjU923BWVv/e384A54E+2YRQOUrZrKSMak3pucoZ+wr
NeqLrDqa7/lIOulybfZwgYeAD0yhWrWuHJafrsqokjm31UmB6ycWwPSFGVVtcL3bZrwEsjCEA8gz
XyWrq97XdU91XsQT6g/XQeLUu5ewTwGGI+wbT7HQ6dGLutnEcMY5RQvGUoTcCcGGVlqUHr4hgn6u
rayTi6+JjXIyZZijoouBBjBaqPRb65zi8GwkzDGC3NFRVFo7PfPu+XLwGSmvCngHzE8pVV3JOqUt
bkAWWg+YNwdvmnxFWdamUJoUDyLaEKl6cjLW9QHe9RrjptEcVvq5DNCHyI/6GaaJCqSkmYGQ49X2
B1UgmfoACf0gXabgBB6ryRel8r/kCa8yegCJRILTejTTDrOIKJVZBIYSQusw8W3ulTYB/zlVzxee
16RfYlJ2KOlpjgleQaOtupUUMClp2H/yRj+jGw9kwNKZqLImi1APA5ISkNMwCBH+MxgA8MUiOZDC
1D6gAaMsWzFuOTkenhLMsLBbz0bZ6TElwgnpqZEEQZ5oHDpSBxVVAwnIlry4tyIanFFAmiTRsy0a
aXDXazCwhP7j+haubX2qZwZ6AYSu5kxJURW3jDIBE+IERtGUgsxFmlx0p4LpkWL5qmnn9Gs6d+fl
COOoDj0RJLB6APvbAPucTHBC1u86bQnG8srM91LcH4Hkex1MNQwUscx9KVUKXDIUmEasZnox7/nz
QQOdHz1FKHdhMERMM4KcmFi0KCq/w/UjPd4crMcrYmygQ49NeMiMzcdkH4/tLvTw5nYcJdUetZoz
yPthJS3sSJ6VvUb/K5J66DEclzDovM9WJuoKWBWOug+r6l9vE5BCXDwFHdj0M1cxsWKPXxcIzu1V
jy/zOfqycW8OCM38zhxadCG1uQKjReD+q31SbW4SVT7s9wRDUN6lzYIzqxMlDDyKtGtLddha7jSB
YInrtY9ZTokaq9jimlIZQJXlDnamo50YvYK6YQYh9V7a4LzaIuCnYMGNKTz2rcz7CNtYlMmuWwr2
g5zqms1DBD4gH0UqNTlvlgAobTAz4Pp4D37ofPLkMlC1I/c5MMtrzMuwSKs7KUdpn5DBVht2tNMn
5rcAR1xNsO1px2cbBS7n28AZwvKYt+xbdqKBasm0HIVbo2vMCQf8c6XBIeML4nmZhFDeFc6bPIJ1
QwbWReK6PSBkPm+NjJoZPXZMPIwOxgMhIHE3NG7ZLF4s8esIPtqVpUO8d+n+rggHV7aptrTTwONW
ZaiopewqtnPuzRyko5ucbDRlYGDF7ZRhbi14ljH+o3OtboUc9KC5KDTvzcJEcsqYl6Se882CA9Wo
k6VTN2NnWstAWAIUtSfxtOKx/O1q4K1drcqVq32HMuFIPHMCnYt7QJhoF5NdHONxECgzHNlIpV6v
UkU9Xf4511DY8uGNVmv10Vda0qn01+bXV0Zap9kEe1RishvLcDdWnlJBoTurwhAQ+zRdA52vVLrk
WLKdeY0gBZLtP4qivQEeBxW9n55r04keVW3AY9kahjeHLQZOHOsDKV3jtAZokp68iT/+Cdgrbt51
GXSVFZP3AuqVrkEbaYtMEvmuC6f2tk4G4t0hjCPnMaxL94VnQmSwfjX0kn0AWyJt8qzwdh14ZCHO
lij7SZnsUAdo0klqPCEoJBRiwg2TcnBwCy5qdBKAK16I8bTt9psT2DhWptNljZ532/vnlWRCh7Ot
06ApGq51bVyUB5YQsEB1G53RZZiq/0YlqML+NI8mtv3XNyOFUgJqF/01kd0/QClhVZGt2bO4X0vu
RA9ON1wWjkZmA+GaLo1oBLG5Tw3mhsAtPdWaSRyzY89uyy6UlMhTunIQu+wT8wdfjoKFmpbGz4b3
O6edzXlsu00dO1JWG7XvrskzNzpEs4RPH6vOn3MfpRT4sT08V30YUcJN3pOJUPXKPPaFhzeocpEw
KGa/ov3+7VyEPAgwR9aurrrKpYhVMKtUNa56jt+7KU94XaagdoL1/iqiryp1vRrAyAT3he9/aJPg
kgQ+bsTvc7Asl7U69xZEZ4VvzBZYWYpEOTFc+4Ul8cQgL4RO76wtnxJkj/zt+pJKbbFHXlo+Ixgm
J/kjfFCR14d8ambg8QC+6y4ZH+ZK3MfmW9d7m6WdXBgwAeSvg35PdZFwBtGn850p5bBaB1KeKeCv
MJTHnP+vzEPjLr2LcvREKa/yQYjXJPsUf/4M40xe4WYi1bRUaWMBvC9kubVSezhXIgZ5tV+SkUXK
VAsFYc82j7Jfyj3MEH7YflT7QHx4ptw9fbkRRd0CvOve5QTGzneSknIACNmXcOOV0RvHpQyV7J41
y4KxkJ21CUtIzjkitmQ004iPDRg/zAK5MvXt0J9VqQXGnXmrz1F22f83czPzMwi8ScYX5Y4huf5t
dRHLL8bcwXNAfBaFSZe92Q5WEskTIaIt5IsEuA6OYjHFQeLko0YApnWU1awMTyO7jAJQXBaRqcC8
sIe/X4/Gb6x7Vw9P0JjeQ6Loe5w9rZoeGT7XQvU+3tNKVq3D1lgLBrDGA9zUtcpfE7V5ZHEQlV4j
u40ql/DQdPM12gjHa6FkKhMyxOMZTr8dHg4SSCuzs3ZraHJmbqe7EROkW36jDTswkRnxRsaU/c+f
HVqoA09ElzzXvS36iPxNTQVe7DfsUJs0S31nRarUysOJ0p5iFPnIIDksCvV8TwOSK1JziV7ftZ8Z
3MCfM0DArDC3o2AlIN8SbRP5PAxGGfeQNtioEqSCOoOnZtqviYHlqETWH6kZfY6/WHDdYXFi0OC3
bijIdo+IFTFyJXEiOtPPYpKpPVWaKTA061t3K3oJ2BxksqR3FrlOui45XnkU8ZbCHulj4S2ReXYi
nw0ns+BeIA8f7VqrPFO4ilx0UuQntrqlCLOGnLDdAp0GD1vkX7hmsYqwr5O3r3rey2xsE/deRW3r
DuW9lwjJVq0mJbxAoFr6XG0P7pLv8QA3Gu9lAG4yfvGG1O4RrprSBRsBC341U1lg4Kjtzv5ggynM
xS8e9Gl+TILgiTOds5c8qtvtiD11ZGgUkjYWXOxrivzWrv+8gWR+YQWeGo1JM5APLRldwUSWx06h
842jmaoq5/XMnO6bJTuAHE7y9joYYW/X7Pw4NhFkgRvqWNWzq5ajnxDviyHkxx0RlACSfQ0gER4C
ZwVaj4GmJCLkKNofzAuHut0hzxv0o2UHSv/z08OAXJ86YU+sKd5KDn6Wj4raZ2sVwt652Fj9CIOB
IcZXcGLc/bQSW0+nYfXgUsQ2WyineFXiCMCrJ/EagdfqsiYrM8w8o0TwebxKk5JouceEaZebQaJ0
KqnHJhorWqap9AMOl28JMZRJgd0kU+g0jdnCDC9D/JqJ25VQb+a5T8Rc4PodPHBzqoaI/Kbxzw+G
gdMTK6UihLlDc30Zk0bZeguyyrAkkdQP/MwnKiZdzNCyfrMVSyzduc/zZd3uyaf37oGs1g+bOBPp
XMs19Y8yvVzZDF6PrvX2RVbyeYZ1C7GtnKXJNGHGH4HWQ7KdjzTuTS3i2lePg246U/OyJj7Sks0k
oorztI1X9i8JBRXc+CgrVtBvbXz4iDTilenDwQcmQDSG5Q+3WCo6DMg6EC/9Qa21j1EKkl9YV7kq
vOqhDgDXs5HVDHmoC7g6H618MmV51tSPxK+Ggx6yoMbDCI9QOKrt7anTD0JMSk9bGjpVt9sEJCWR
koYV5ngYQolMD/t6ty7UzP1BwJf0Wfa5lKU5dpcVXfHlUHvYPWSVzFug5Kz5NPE4qWmyIlsGNZT8
zYNxRUjxz0/4hzqijr2r7MG1wx6ABJkv72lcwgMCORQtivm56E12f1UM6h/+Hw6yc5ONWqL1oGJM
fhfZVYnQ1OaX1GNt5zwlKybNjSBhrE57wghRnsb/WlsJVwp7ejvfyDuB519vuABaX9HiHbQY+n9h
Wo2fBUcZPsKOBKVCOAl/S+Gr13DFmIIxxh4l5AwrRXi0gS5fulhrSl76egqcp0cRbjmoiJOqItmz
m3UcEioazEhzFnw2vMBVMlztFwlwegTskT664UqLb+Q33C2/x4t2eWMEUUA/9rO7JaP7E2qaP8WB
LbTu5htAyRk85qxiJc7B9hO7JnmBF7ciVgZHvMIASFyiT1BPtVj1kSBRmeH+AeasCR0ygs4/L6aX
kHRXicqJElvYNxauJlyLC6HpIoMByLDEEMddMrW+c9GBxWVjwDbAw9fX4MM6lYQMZvST+YR6JiBP
JbYgUbQyK7b+q2uuwBGd17cIOXztdKWurTYCcM31yZMi/LHcN8zjHAd2aPhAJUB7nSzgEokEOUWT
+RTgqxiueT4P66m1Ttd6M24XIrh3NSz5Ij18SRO1J6n9mppZq+LlZ03gBswRbRSaX9esIFE8Pq0N
z7NDBUcWZkf6KoKuUPFjs0ScOfogdJyZ0XYqPLWsweKx2ggFeRqpWMUujl7BWMc3K+VkTB81sAyl
Llz9DNHToCx94OIcTly6L9GdNjzAU+4PWK8eb6zUo7WvXV+a9UNOFopmSNPrtst3DGuVM66Orj4x
F8dCUf+qH9eDHhmvdTpGnWwgjQS0+3F+70fGPJNhkdCx8xftwhLz3Y4CYEFPS5rgQoPh6kX53U7k
AlIYPU1wakQCirFbu1Fcr9Uz/BGTsAK2E2TBpVgJZPV0Ezpl0ifV16jk1hMsZcVkcKoeY3Lw64SL
w2mlIUTltJv7MXAH2GDeBZ3hnF99QSfOo20fzimEd5TzLyccFJkcsc679YHqP61GotVEBaQ1potn
iCfjPWRoPz9w6MYaxLEtuW73T83yV7InYedMdgU1I9D4IaZTN0MvjMck0R0Emmq4ql3le8qMvipf
vA81HXsmsOKfJEL8WeXbD6XEqyoyr59G2Ai3VjglaBtynCwxSPWA1/F4W65Y7h4Zb9+3CWIFNOdA
k0J6lG9h3VSwt1aHMgpaOdPV9vrkVBMN+pkMiEDOvnbVqJ+CMd3OPLEsh9oZe6C9jNivwMmrf8mG
2WNnLQ3MutW0WzBnQNp3WRnJigk1fMJ/fmpRq2mO9heIred4rIJFt9nP5UZekAn6RgAqRzNTtv84
XWN5H2eMtphKqRI68AYDe8HcelEFVD1WEOFHvfVJL9WZCfwWWNWtVVkcnVQVc06WmcDpAfgnyLIs
sy3cljDjCIPsyufMQQ280j06bmG4gikjaSb8l6p+yeZk/PA6xVxZnXmYfzkpKPAnlxNIqG9/maW3
eHZT07wJC06podNlhDAqpCFMl8ns50xC4QNh1RsCxTgDfoQXC+o/54hbJmv2ahrj6mumu9dxtbAT
ikbMqc7UUIydtU06vBfLfDFdK/rHudptwsTtnEXgQ+4TqY+YyE+pKTRuFPohse/ySCoFXRm2Fn1l
3X4W438pY0cOMHvsw00g0CoX4B0eD60asobu6tSKeoxXRzp88bjfT/R7oaad65GPHL1oeOjMYGmd
9o+FiAK9aUjRUq2VWiN7p6cpWRI82Ugbszz/blBmy+wWlE1F7ilOdsGj0gj1mza/vhl7raAKO72W
TPXA18in2qNHif5J28HSMbqxKgrJs6GBqvhdLJWFXclNVLJXed49BjagK3AITRWMqzUDzfDgE1UO
xv/mjUSCLu9ucUzZmAPOqWtaDjWR0wxnK8xKncdnr4htfOJ7pZDzW9RcVkfwngsgFbEvUXj3svaZ
U6RNn5FaB2LcX3LEQ14l/sYrMMoaJXtC4AMsZ4xWKiZ6wfMb0NE/9nnf2qku44huCisTWiURFPCU
ZrAme3TCRuOzKMjSGjMmZHUtY3/CSqX3zSHXmqDjuNhj9dZxAf8kBwUWGpALDobKSsAgOc8Sb4r5
qHCstTBAtRGdxhNjG+n2e5hjPF3T2KEfipoEgbUuzZ3qysw7JUGnZsdTWK4aOMgoVfy3St07Cp/J
lGyAZMcCuHZfAWK1uohMZbwp8ketgYrzRIVIP6u/Ynl21n266oKOftA0BvIF9Vzl1W6NH898N2Gs
YdgPz9QmMOaXWYOjTqEJARo97LIVJujf4wbKwvrhwq6wC8uGDEwuScPRv/RvNlbCCegrNF5V3tb/
KTbglVzpCzCq9DtFDJUTFP26Co4ZCCwgTCJ0GJAykqWNgc/YZYj5ezHLFVCIv/yozCyH4iTa0Y10
yQGKTkGmrOoltiaTCaZg0L+gAOHHf9zEIrQJZm8v4vBuj+B0RIhnUvKnWka756IZLvejpUQVaPL3
5/vBUeYhZyLYdyHxE4+8Gb5JA+3rdOZy67DmvZKkZo6+2MRj6MPVIiXd6Fl7Pjz1Zr31hNMiK8Qr
loD9YJVVx0xnxo2zf4vbjgec5zbkpDiWtBwY958crJ+HXezCqdEvhuLggJNSDljyxiEyNMj81jK1
tGoYoMfakwhun7D5VsQQ/WYbpyekDc8My42ordGkKoufIhGnbLDubyX0+hIeymmDANM1Pi4BwCOT
KgS9DnWfo5h71Tj4/JtoBtzT+WwTXesZULx5dNnyuZTk15akof0HfiDCyNEwZbFvmgFW9ZNSaZKK
/pkSj068KCg76lZZTG1kTq5gA9NUbtZuSd2y8FQbTj8GmcJSE72epgwR9Ialesb+lEEdYmc+krSa
RgO5EmpfNPaYEDwvYPLs54Nlp68bVvyx+4hySYUEkyyW29+pd3pigezJ9cr4PiqJ2Wd0tZ3IHfax
N9jboVXDHSajeMMgiKwRx6tUumUbArkYlCzTflJnAPCHCHeJ6DqsuOZnVp+wScCh+J6F3bBmrw1G
KJCDHRgdW423m/k9CjplkQtTJ9TTLTEa5Jnnwt2je3joloUHPn5dr8FaQMP8B6wm/hr0BVPEj3xf
QLZA1ZR33YeAN5NQE3h7CSE7zb7s65PyYgQ8qdyx394x4BwR7B8ymVcpLqM6K98w8vxBhVrTNeFd
e0rP2p+8lHMdo5+tA/SWTmj5chr07Y1/vlSURsZQKxtQ1OublrVE4Tuu2l+Rm4FiZEN9ZajLNMir
c92nOhBfvWNN9tySo526+FDQBHjD9V/SkjNtChYemrWbq2/CCeuleIhPCXZrHQQLtBAYrpod7GTD
wsyWu2ZmKuUvsVk26pKvZq92zHWz58JYusgPhCpb84Z+rSlXW/5Np/YJ2isqr2VsbvMN1iBsUqUl
Qzz3Zaxp2W/r5Yrgyt3gTLawUPB14pxk+mRI0ZaFQMtJ4s1xuDRvjUbka4s/gV+JYuM01qINSCbt
kJD6pybH/98kGZg1/aSu5BgcCeMovtV30a61Z1H4gAi+JUZk/orotwtB7KfCtfHlUXNpdbQxAgyt
DFA9YH3f98lCgMgh0D/7R75ZDWzdlt+TybELgC4k3BoTahhYJViBbQ+byZ1vW02NMivFOhYpSfMc
mWsz1Bt18aGCHazJ9gc28q225ndq/H5QDHKbVvNJBOZJI6UBKC3difOrK6RQO6Sl58Y0+/ifufCL
YCyYY6uYgqqdTmGmAwaTuLvI+HstnyCo6UmqL/8+PGDpdfNtf+j0PD+bih7SXRPsXBaiD38H0QUR
eHBq8NAMC3CGb3jPbein6fJL/1DW4MhKNOFWnC9Y7MyqIVnbD2JIgQORpOtWRuNDZVB2iwpYIj+Q
EyYll2plIr59pcv+eEOkxUYdDPvjE+ye7p61b/9SM5A65XNeFM0gcQjxN8TpYBxSK9jtRa5jWCO/
0kmg8TmZU7fYTDn93MJhNHx9NVogGvRixj46OXI37jwIDI063yTnYGN0ARaDwIzqHnISW6OwBkoF
a3WtBMTEPs4fTogiYgGm3y/f8a87jn4HDV/jiz+1gDhMD9+ewjv/LEzZE5yWOoSwMVyD2TNtY/vU
+YgGCDvBSHYCxGwSl0ehrlbkVsyg4XP1He5JcNZRk9OCVoxZFcH3609zkPSjTeGDF31d4Hdg9dZv
wVC7lMxrTSFKga6ROeeITsvF9hu5Yxvo3XLvVx5TdkT5ILVFcKFG89WbiRZzN/dsJxoi4+NEL3hF
d2ERJb+f0IzNYdcDZb9x1pbK5wRQheyTaGt9aUycpDLDgJuk+Tmz8UNpOdh4yoFPjg2/y+6AxgyR
pRMt3Vnjy/RY491vQzAD+0C5RCHkJFJ0o6N9Wuw54GKMfDu5jhpeGk5gR19HwHoXO+Fd6AGzTNpc
cCEhzkTCKJT/3PBKMUZfz3gO8pdfsrisxN1QcBPUUnGjY5Y4tMuOPeCDM4DeK5WaK3DKN6Xfmk1F
69vbvC2d3YuIRkLzaNSGekCRk2fM8jQ3KRszrp89JtDkvZzdzh5UEzPYMWUzGKi3geI0ut8uFmpW
Wxdz1n1QvJ46hNryOfEM9dPTyalTK1EiUAQBN7yWlMHyyPJUmt92x5TWJ8+3iHGRc6WACMQF67yg
L0iVCqQqLbah4VyM+uekRELvFOOxla3ExY/h1vI66aVz3d+B8MrT/J3Xt26opRSMCriLyuP7XgTB
UJ2XlEbdR//LjR17d0uxEonBWOx0opL4gf1uEJzdK6cnLKAfWzu2uMNI58wTrLqBiGJP6S1RgFtr
dUBPFZUmN1VtcFU3JBXhoSAL29td57FPmVHTw8bhGc8yiQOtVKnJrGc0ja8ZRCJEAvxUItycI+av
4NQ9UAElc90/Prj9FTXFWpz9wAJCSkAAFKRhzLvOdoRJ7QNet5cDy2oAqP7uKbFdpMxjs7IrZ69o
shrevoSoCTBysJqswMEAmNdaWbZ2RR7LMTsVZfXZ2m1EQLWE6QVES8sS0cAOra9VwAXN5/CMJTWz
UZ2u7kbMFSftzioYyRw8QhU5CFdDRKYGdQv0r3o3V/Hg3ic90SsdT0x/lL5BjypiASGYudBOQcki
0ISX8Vbo1e9LDG1PFyPVO6TWAypQdq+edEIYqinjaf/YGO/6GgdvxvsKcBK6EZpD/NM0VlEby3Pi
2bDnMSg5SxfM1akQNqs/Q7KcFiTLQGIjMf62cHDSUmCRzlGHtZAvGMHyU8ISDi2AutQdpLWRvcUm
OcOmxewQ+Pa1jOEqYs2OOYgmCpAACfoIdV29uVYHi2Ongsx1ftkWIln58/L4P7TNby6ielZ42yz5
l714fROMhTJq39m8/IXQ9I6bbBUyFdB9OhUoeym3QXSfW1FT86UnfJK1rSX6HxJSHBb2Cku/qhmK
c5pHgSw1qUYHmskoL9u/ZZRdEmnaElepGPolQJ5uGxeQB5Nni+6x0ZjqDUSUMCWWKzEvELOzkAa8
u2W9MLQ2TjQVZcXvx/6Zn6tADS4omJJG1IuJRxdKo7X5PaMtrGRGs1nl7fJ6fccmLkVlspvZsSFh
cq9ApDDSl4ZSWoUT+DRC4VsYcTvyfMxaGLx3PvgOOjMRYuP2WgGQxMCPbhJi4Wz6UwHMqaN3lzEu
gdNMLGUCZEGUP6hecHK9O4uBP6RkYfTkO31xkTJuq1aMeH/QJa3TjhEGB9q9rmr3YLYpH6he0DBq
Kj66J0iqqd4qpbcGsfcI07l/5FnMp4RBN4JcwfPLChCxR4Wf/WG5tcXU4BjtdeGHnLymctmOv3vP
me7WbL5RxAigxQHKN1/9j0hbZiG606vmtW2zQ3VGQQPEe7tt4PVesARBaiSC5Ffih9Q1LVDSmqlB
7DwzpP0knEbqRUHKqlRv5Rm1azyI/B/dE9qE02jDAyKxJs5uuxRPkj3TbhAXlx3r2Iba7/VNiAfq
Ct8nfA4pR3dlhaF56JYjjMa05Or6bUyuT+tZGmzyhlo43Sml5JcoagC32bF8mz7BfyrVtLiSWFcP
95iXBgRouk9+c6bDcogYf6p9W//g1aE32Zt6fOf9jc4W9HXJWcwHOIb9E9emPWt2aeZo4j2mf+fv
XFzHlUy9YjKBQJUrkTR4QJ+QXfqmxTS50O4lrhipmTQw2flrDgXZ20sNQfUxmTkZ4tMD3XfqiMUo
gdz6v3qEQngBkoKhbwgQdKogcsRA1nfSQk0rrQJR0qu3l8N/vVme2IxhXo8pR5aJStT+O4HUDf/C
w8/BV7SRe9DqJmXkrk9EGd8laXHK4SLHWCNdKjgZ5cHr8NBIlyClouTnkJltTTCQ9eQHA9gAszCQ
Q8zzISS41nT5ASdmr57LLjZ3gQeDbL+ffh0cb7wfW41wjL4dwTz0Ml2UG/p2C7C4Z8snHahBs5sA
iFUVJpQfANc/BGrEQM+hN8o3iNqtHpvoKM8qljEryrRyjjonI15ZSrahkR9eMjg3Uk4FWspLPcqu
a/XYO8A4YNAxfrGgKNMkY9Uk5dEG8HzanLI6vx1pQK3sD2DVrXt90+gfVr1WtP3lZAhctPgEHZfu
D3zpkxTCMNaFJvohpfXH6Ko5nM75UvMdhxfa4WhOmspFkwTECkZSt8UpX6/BiDqdZh5ekR05tgYg
RuN0c1euYyT3Lb2vZUpFo1mXTgtL7qsyO5FQkAr4zUVzaWb+nEOaPF7iMuPSLt1PCHXycxpS9FHj
eRaK7kIO1ZygzKhAKXg2PwBtoseu/Y1N4NX8CiDyQZnPpd+3bqHCXtYK29cp2OsrjmLiOAI+AsPW
MEsm/ij7q/TnWL86S3NriPv0T+R4zcLMepvYsUaf3GwsRrRKZEo/d8iYj7DhojwNvqIak23KsPtx
89axYzclHGhbCA2qjTzLhemgB5zDlqriwXbEQ26LeaNEgQCOQkahxIHdkPU23bE0LU16d5cS8N4n
5aybW5rbXiSlisJL28W+PJeKtBuTJk3zcZvlc8Zkv/vkojvzNZDNEoPbJ4T0GKQsz2Ejk9LzMQ6F
7DrpatNJ1Z8DQYLJ+YVherF0ohzahc+q63k6kGRNBk72sUuGFFnLXuCVL3tJQFcYKZYI442n65hz
LKO9Xf9XBwYRURzg2eMWuRxElKFS6coRgV+ax3flwNzvFPlGEWMq1+7Lk1+M+9mRwlN/B13HrzdH
lX594YJtYBPm4KNvVAd6Gkma5Od7QNgf3Gd6PO7skzwXE8YR1L9OAwRcq/Mvnc7jW71i76svkrNi
5xz7I10vIre0ZL386QhaOdgH3WX/cAYT1vVKvkLHNGCeQtterpRl6nZhg7OHHjuBdb+BUfB5M+vO
3JhXAxrA+qeollWh5qQ3RdM6VVN64BEAwlKqmSrehZLmEBksWoSpPzvlJE4tPhDbXr/E42R6rlef
TrwlmPoCJ6mIzWAep9GbYIyjXXa1ZdHKWBKXqjKTLivvhL/ich4OMS0CHH0WdbSvHTK2ZAEpGcdg
78R/i1nWY+rcK4zOFuAH0MY9r6DvuuflvCDovE7N7aBsaY7q8NUMNwGvFyxai5IZoAMuHgLkH7Kq
2MNOdQYY2lHmP3aCiwQdPF0AqTwLpz1IIx2golqIRlYhmLVlsy2XB58BJWlzE9X1YH68ftl3GP7d
ncAFudx6teNvTdjrnOb/7m6TmMVWIwlQxNoFfuXGpJQAWsso0xyCX89MQ6uldscnbaDIVWRaIAQX
PD5DX4EtjtVQ/nKDeoT7gL4B/JJ5aAcIehxz04IizW1LDhEH7qagOWxq+7RsE8/DXjO/XR68+SMv
KQjuPT53tFh8ai59FycMXhqTALbb1REmsENaKPYiK768ObaJyuQLJVGXqV4zDH53SSWfcOaAB3pB
sXIVgeKSlrJTWcmuk9naUC5+LXDzspEnh+uPIyEj8sU+ySvifbwYgnyoCkOlnek8O8E+Bi92n9Ax
WQVWvV++ATDMmHKZSWfNOqnMx2S0qj01ct5rTm9L5WALoGDJS8GILDPtevtImR7WmsufQ829hG4S
zZV3Ro2Co9Ayld6YXgInw/wSwS14u49wTLxTJQ5RiwcK19jygl1PirTi45Rq38bwiKXS0BAUXJSG
5jiURd2yfSh173V3CI8evT6J30ejZrGkpzUZ5nvGoY1Y+C6jxjXESL72cf5qZnIUiA8VUFHxVh+p
vP7zK+78jRDdrFntO26pjSmrJsDTLNrwzsbcKpnFVpReaOn6wDD3IoQOPE6OFIh2a/0T9m1R1r+1
bLaS1c6LPhROpDXW35d6OcCsmzMUsL0Dm2KWi4bs7RtH2hA/hYTh3D209chlWbRMSGxszRTJ+z62
j4vZABIUNAk1vwDs67NZkPykc+8jGAI46oAbZ8a+EefStuqOFlsWTBXuHqxSiKFFITDXI8iKKSgD
mRQbaC17g5I7LF3ISonQoQ7lpjf6WsqNUGJDmF+fpJqgY6U2QfNwYMdBwiq+raXseHZRlGmBEIqJ
xWRAb3yddBWZYBw+qhMno2kIDOSwIq/QMxEb496taRtWyfA9UBOGzqz6Wt/RhoQZNms+VTZbPiAT
B++VtgRIdIo=
`protect end_protected
