-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Dnnd9AeS4g2owjFXZVy7UUaNZ8mYkNqcFseZhny4C3JCcqSYoFqUfBpORHEYs4R9EqL2ZSRq1vBF
DZJbIeYmtLKzTduJ6s2waY9PdTco1kjj3Vngp3ZpLmdvpmNLEcglIVOx2BI4G5ekUn0VRKEGPS+W
RsKI8jx7SiPsVDd/y6g++KsVIaPEopwvnS+/mv4ZbgS/TcJHJINDfbTh5KayhJ6K43/oM4GWkycj
smv8vzY1JRWUcq+NvTgW8zy5GE0+g5jO9vLBJ9OCr3aFjodvZvBg+yhzLjUspnYvxWo29qHDpKdG
a2YjYQAVCb/c12ltHMOb4eiinb4ZroyWKBHW2g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28512)
`protect data_block
4WhJg68FT6rxlc7zR4sTOG33jo1PrijUgzjX4efTudZx/KrRNa3EU7YS1UQVBfB9qi3bjbJDGtS5
zW/iybWCK91XwKlDWNmGj+InMuv4AKQDNl8F7h8JaUQ1ZL5jlQbNZYRUieOmYCRt+egWqr8PN5u8
MCXAwM+UBaQ+U+WyTI41+WcrddKuzpV3Qpnhf/F+TN56JFnWQba+4ETDajPjwalZGLhATjKjNHy/
ZGjmMqJv1i5OP623RkMtZn00WmDlpdwc1kjru1hJ9d6JMJPJpv+ytIly2Fra48SrmJGMMrOS6wLF
MiZ5IeVS30rC/VXCF5tRfrW8mPpI/db4Wt3SJH2VjSh363iPxP+1Y/+bozC6cAgQyfh04al9a/E6
XDMC1Uygnf6rAfu4/KdVXseP2kE3jqm1CeqbNBZMruor5B4juoTTLhvXtsWbQoquERGLn0y86Wxu
uRtlTS2clNrUCalEqLE7NyFgz0uOvt+djIqtMme1IUdIfx03cyObE5F6utXESJ8NsEPti7tPxrFu
fat/WeLh0HX+daYPum3lPSjCnaP55xEu5RQABAWBeRGlyzTtKOBErgT+osQwroURqDc0re/dME0g
URWk2cLUoHwiFk8rCXK6wlCGHbVgXQ+jO+yp2sYZLSRB1aa84zrbCd/aF07xdfbu5q3MJpNsBB6F
IilsKNbQrCXhw1hJJ4l7tmhUYVJwd5Gz1BQ6foB67lEUMMOdXNGavvn11qVhULfp03BElmV+QPpw
kHyW/HbB2Q18voIrKVbBfoLltMZ1/6AOILiOVw1E7FPvAD9Gy0A3QkJVfNE2wp2lEM0lf4b4ULkv
mGDiC9AoQFD4i+lvzIV0WMxJsmchcIySQ/i9AZYUatwJ+4dBgZc4zUthtj36L6vqreVHAusJhe08
a2PJ8PpXb03kgipaEUZOgLQ4Up3x/3uZoac33vhPg8yeLBj9QUDExVa8socLrYf3YwEA+y6u3I7z
VtqQAXb+U4rd36/w+IYkQU0j7JuzDIX7S67sS27Hii+hbRDZzJH1Z3Vt3OM6TtSZ81Qk/Lel0jWx
VGyZzjCuT53JByH7OEpFrJIxvlIp+O89KMcJLP/IUlrgkNANakFQWzZ3MVFdI0y9oVhK/2jDs8yH
W2FFf6sE0voAL74jhv8uqJ6WfMcOQn8OtqnwYzjJJtwOfxrLm22lqvJfIqfjf/KT7teQDHGAB/e6
+VZKp0tA/wexyUbwDwLp5Df18G7nO/qc1BeBVoAyPuSu072Z3Qo+dDSCOEJPQ42Bm115ajUzBtaB
eWXjV1c9yTFRdv3k/e3sbfsRmjJtecqOQ8kBgH+9a78J3Lop/7QZZUJV1Q5YlG4RWrp5bTWwP5kI
/IAt3vmFNqaBUp/LMRZgZMW58cdvH/0uvKnuf/GEB+WtY0VmI9PiZyNdMv+zM8eET05VgW7+Hn4E
BNC3dJXQn20ZG1AJQ+W8XLL4teGOLpY/1B2QkaMuBiN4SQCU9gzju4JNislfy7XT6nmZOXSQjjGH
9PNXcgMfGXEAkbzaB4wzTAVLht1nAica+/X/obl3DB3SWZJtIM6RQ8keib+sa6ow22OghkS18+xv
VHmm7lc0HaCUn7dVahQYmZBhNTx1H+z89y+9VaNqtZmkB22u+46ogkGfBPcER+Do1H3PaqzVZqNc
NrKfFFgFYmGNwGfX1GY+mDLfERst3O9RtN0/t9bdFLjEWjgUvyOaGvCLh0pf1k4AOsjzaQ01ld8J
9y5DrRAeUCxgRMoQY8rId6q53ciYcDtaWFHe1V+d0uuyDB3TxC7Tg30ZovxUt7hZbB7zXo+15l9s
uDG476uaJDAN3pKA+4er5C8f5KgcF4SXXkJB0EVG0UUCDP/VoNCFOIoBYqWJXIIM12zPe7I5flBy
U2TtVgrW78K9wr3KDVA0QACD67OlAHqq/c2LyPF0gQH7/AqHpKyuNSwD9ZztlDuG4MrCtcylDdGM
nJmjJtufnR7y5SZGZGuxuuFzAcl8/r5gP5F42FO/vjWHT5lS2FSRH0ojZWC7IMmcKeaaPALrEja4
34ICIBWtKL3Y6VqOjeCUNEmon3/ddj80RuxcmUDb8q19zJGay4StnWKsH7Us6dK9zyDq3H37ra19
EiOjw6yJIEUYsHcBW277+dhmKsk2wEqqxu+Ew+zcHtxbv1T8fSNeSNrtVstLPQWosDq62SbaQmBG
W2IfVUO9uxg16oy0lJsvlpIKRXA+iEL8ipPr62kkPmEQWoyy4Epe8x7z7IqoFJd1GGg5e4/CRPm4
OvlvRkzkDRI1nFbOnHQXN3B7BsAC3i5E8o4SkOqq29zmy0J/HVEVIOF39eCLBvoW7QVxfC2zfIHL
/+Yp+19wAVHzq4x0SWGh/rZ5wpjP9k9+lH3zPpYV4CV3CdGpb225S5ovi7oj8nvc0pFCKmc7wt+9
HLHh+TH44QGyz5lRie7q+uazXc9cd0dAiVMDrk0xuiZUaPJZ23DwxOSm4pTfgJ9pLqHkaPk+GrHK
e8+syqq+9p5nVWMLHjNywXkEPxVvLp2ysrKjIBZ/NaGlYaVBtjCC+7NdseZ5ZhZvyPragb6GwBlw
Mz3QVUR9KuuuKPInS1k+I2vfajBLoL0c07LrZhS7IIs5fcj4VzXrIs5POnl/8iX/fWvc1akgqLm4
e7x9v3iVGFlHIpHtxl6by5IDaPTiLwkkx588aR/Flt+guXpZNMCfXK3Soq8epCfKjguMrhZDxZr8
m9lasqJU/wawhxiEF3IpyAhE8brewTLB8wtsS4CDsdoiy/xrWaWcTqgxr2Ku4kuLKM3qO9Njg3HO
Shmr2uFog45gIgjQR6EFUxrnhcn5OoIn8FZCkc4BIuKayMdh2j9ZZHDMFUeFEs+GsAJyFzkWWs5E
I9d6zAI0HiA89tDXMLSWMd5nbfc9UUPRAA01S0R0RiC132uKmO/t8jjd0beHKssY6hUBb+NFACF/
b3nSOtRnbmtJ/2h3S96cLj4g7xtTPTswx3NBn15MBBVhNHmoaYqULMtGaJOsnQtIpQ+QqyUkooIq
Mn4RME6CM33uVbqebUsLvlvUjsyPtIDWLsAoeHNGzMf/vMgR1onqfX6/BpWE0b4u9jjckDSUWo+7
yaSYKDcvRUaYC3OSF/d52CG7qWSUfnzROJrLZKzSpQphL9MuzE+cKweQ2CJdzl/YYyU1Y1b8XU16
siMLLahkPJtRg6u2OycI/oAChum0CPE8+qwNdMfHAXZYxYq6DXe0SDax2EHvRipkxlKBKjnj6JPV
cezDDTRaIasjrkh3E33kGB0XmN5uCOF3tKfr1dqaiPuMoFSt9455+/XwLkhduudK7oyKIBtNgAf4
LV7Ke5etFYMREuYuafZRW3w3dYcyS5P5BilJ7Ah7B0FyNqyuLkJSUzZAaIHAg7VekoXdxa0aoqeW
/GLexvkrdKi2MdHkEOOMCBaqWCVMxPgnD3UkioXs89EqoXDY+i8WlFvGGiVXShGlhO5sdQmtgeXY
DDJCrfe/BtinfuRdrIhavzn2PAVrIPteP4vU+8xlF60vO22Gtp/1+Kdw1zgoBqofxOwRHLG0gbPb
qKuOmiuOWVpiQ9q7OnrcnuekiFcrQBIDBo2knWS55OBDYYInFL/ijhftRHftZ4s66UqNviilkNCa
+i0NIc70vKEMNGiqhUOmAukK21nfjjKGqtwniM/y4MpYeGgLOp03HTQPRR2J5df9lTOzM/twjpDx
8Wv2oZPdf1++iBCZjTUq7uKGta+WEldujXXhB9pKac7Wia6j5nztMA8/jNPovuGsCZ7PAE1U0gzQ
MFtlY82RlLtx6lDnNbzN7QzuQlURH7RamttMRqsKDnnGi0q/nFYwnodwhKcFBEWzaUYamH+rm4yK
H0Mxua/1fnobvBy0lzGKViTxrzsP9fIa94+ZMa/kqSfUFOsYB3fOaBGvcfLJ23iDifHIau/nUqHu
n+8qgroMv8sJ3tBPdInktrt202r6owviFA5Rpn/qnOUqGSD9EJT7ZcIxQYUvx6LLWsQEuAKtbMWk
/sKkGM9ixrDIDd7M/n+excjkjHw6dgtULdJYJTIJ6JUrNTPujZIv2LG45SjTolwO5Ebrr7WdyKW5
R7gnYKidgRoP6fCBJ6Fwt4ZnVVizQbXVhPRVJMb7GGwEwBPJYU080iB30i9fQity17ticQcIQLer
TvJNTCsI4eC1egQCprJ6J5oYJvB3OK/57Dlf85AQlhgGgkMLrRJzmvXTxtKKgMh4vojNTk3exB9I
r25UrcnmyjxgbDGQ/PjLrwhYG4zQCs+Zs2zU7rslp+34FeJ/cNw2cqYuT7PhfJJ13P2A69ICHv5p
QKozgGWqAMAN3wX/paYo9f/cuIynIto4O8eAl48isvxN1X+x/aF88yQszxv4kNa8TMFmtz4NTJV6
a6l9BbEASUMCoQyt++pmrZX49jQ0cVsS/f9JEpg4PZlupBSM8dGrGvXXWF8WUsUwpVHxO83xCiQZ
r38kd7MGsf9VmmJHi+91FLH3/Pz8LWkdvf8hF40C3CgBQ/YDbqfdhJ3fjMs21GD3qFNvlbbZwjuN
uNceaGiUnHxXeD7HZRet+IRwhWXn/4+QLTONQsQveNso6P3ib9/jtu7I4quFdxREkYasGbbqfyi+
LWC9yU21acURhXuW1DG3HbLljqcay/IkIiSwOzDBXebJnE6T6VmlrfeAoQcV0/4vLf9CPmfsBt9d
zQ+x3TPvDVIfUnRhuNZMjFwzU7Ijgr9E9sK/BNYdKRo5fOJikQ7zTg+jCMv5SfFviINJopGhbN1o
aa3n0VQP5aCA95izGQupB5PZYt28SWgoopCW4sTFqQ8GFCUzHB3MtK9McAvYzHSkSQn+Az7hlvNI
PMKwf44vwc6R79ly5H7nU4F15Wz3E9QFdaCecHWznAlojiBJvSgh6sVRSZKJ1dwvREVit/Fp5sLH
Xys9SBbdZJkyvsiXTixy2x+3CgPfsoS7092EB8JvQG6kFiASR/rn1TW/h/pz87e/BDh0T9EUDrFo
jv6Q/5I7Nt9rb03Nl7v60teD5yOZtNckGKn96Yslr/HHtGof87bHNYDrLnqVTTTPszElMUTZoTtB
GC9UJ8J+Fi2QJ+cpi1juwPk6H0dQwChcciW2XSn8XtlSmR091NfvmksDLgV+NRyw1v4AIdsl+ItK
MAb0gbSXTUevVsOYJJGJADaoTsmI0i7X6OtFjQYrxKqT4DDiwPVrphkqFyOiaTSprt+VmR5GUH0y
gQz9xWi8w/RSr6nXuGIHxSChtxc4r867RqSBiBUxhXjZLIAf3F+/ErYBFYQMHmsTNIoEvE79vucS
1chlu/Wbo2De7A0S9Cbj7aSz4eP7u/wYCqH7nqy4UqM84Qadb2k7jVGu9H4NpGqSXHreJGsVgWKe
rz8SmRtiZMe8o2iKE3DJ7SDgV6wTejCy5Rd7vImgWairgOj85gGlol87I86zY+ytLUik8rX8DpGY
JZFDzk8Ofzk5iWYMFwjqDu1+uU+SAlQYCh/lJ6Jhh9ZjcKi2gjZrWVhkwHHf9YTYbrKjfyTkS5Jr
pOYGOjMVS9N1kK0LlhIyzN8ONi/cigS1++cYC4b22igvpvPIweFZ20oZ5m5B4zu9TQGwUKYjxG1i
r3XGLQywT4ROJ2VHiXfjpE/5G1TZdUw0BKLNVHLmY32KtubuZ+9r8554CWOt0ARlC7Mxr6xRLscF
BlbXy7MPAdN2qVHLfD6IPQ/Z1B+EqzSSA6rwFzxbfl0uThhr+KzG2kpHaXjb5aYf/fY1sm/PZpnJ
l/xBJkru0N0etMOCzwBDpPttLTAYMopRbOlUqLl/2BItzIpg1vp1AZsrOmUXUbHQZx204eu82uTo
N07i3qqXzKQdsLtGC3qlGkAjU0uB3UeCU6mki0MAcASJNfdrIKwuCWPC5s34FI0Rzvxb8IOIhN34
lEkz4WEHA42erOj4wz0sDbqDAWJGHYtqV69SDi3oCXvLzVFTCuowuaQ9KLfl9O+xVa6WD6MZmsR/
bLFMwLoIPloO6KYJ11Lp4vUzyONIs65wYMa/dzPvgBwkU9FLjglVqyyljSUNUrPLuqM8yVKgv32J
4pF7HHmeLx5oJ/BR3YWMREEwEz92BBFYpRuDiTAi4YHgyvytNsBNAYWweZKGegLyVQiF9WJISA/W
caMhxTH+PM4SA36YxQRIJmQeDATo2oM0P8vXbMIWhYrdQjyLsW/pMi24C2tDH2ofj2G53ELyKlnL
mjr0A0sM1da8GnSoJD5aNQPX/ZG5sU0XJpNF846Y80/fPBXKmnFxuA+pxU2HWh5oPIousxmTc/Mm
xTFSW3LmaVkC12eeV+eOWlZ/k5MvX6Znt2c1n96M3NyLZWguyb5c4qTnTzTF5AvFDc3GGQZryZRC
x21eZlqPB6qTduQVcDzXu8/hYGtqsZAVy7cJajVyML9alQtNYPaXekT32ov+NivbFtRIvCTc9ZJ6
JGpNnSP1F24zx+6e9J6XQgKu2U+GSWE8w13yrR32xEyRqweddJ4xQ0esZ7tAFebsUxkOtKLxhSi4
wlqNcsC/m1j19v020MozlQthDkLswyxXRf+1AWtJbjP99aoyhYmDKLme2URWC/t1QcySFTkmTgcY
dzFPxueaBDP1O8GMlFnV6O0qwycmk7ejvm7GvUXpUhNnQciIPBXEhREGoqaSpSReXRToUB32jEhH
FZY50EM4ysCrRoIbK4ypwI1hS7K+RBzMpZI+u9YlLflbj44eQJm1CNVRhmm/Bs7RNsKWfjP7/NhB
YGDZIS8aio4e1WcQtqONSrp3dT8N8G8LBjYdD2ZhGzt++3KT244lennIB+kjdfE8ElUzrzVUuISs
wR40iE8Kp21HzYjUfu9olcjJ6n/LHYHMiWQZb1zda4XqoSx6VdDmMmnTXD3mu0cya1E3xQOd+Cni
P0LUflgO6Tf9pd+zrvVFrWDpKxBU9bUUG+z40wHJsYYEBxYqcdgTqQvJL9FfiYBU0l4hiHVbAZKj
j0iBg/uTJ5wrMGMvuoDgtq6UHi3k3QeSfRQXSVIwy45uJSpyOdE4cw+7HqfL5rMZ5wJnPIwwQtA/
Hu/GvNPcYPFoLhdx5DP5cuAxt1YP/PnTYw/777ZMlxHgTipfFtj4YHfo9WPNnFGB1Z93VIZy3GSA
5O0zMvVAOKQAX7otgbPyoHTiQXhg18iOLR2BZ4DYw40DvDk1aABSWuWts5RUl/jd3cCTnLtfYUHo
cxwXplbOCP0G3maM0DKIGOWKJlyMBU3QsAkiEx03K/4ixaD4w0hsecXTzhwH2X2dPFIYasOQKAm8
JF5oKcubuFP3Atn/ZXFVGi5Dt33zAQdOWp3OQ11wH2SRcLNfc6PgDC+YS8+TfvkurVI5DUOihiod
WSRNbYSNTtYMP6H6sZ8ZWtxaADXLqRI/GHehQwoq9AOtxa1tg2SWF/qCuj3cfKUwyvL1+ubCfuG3
Yp/KtLimT7nmKQT4lZwsq3Z6XIsWYPbrSxIyT7lkl4mrOYpM2G8KdIZlkQ099w0ZoGOnfcyslsgS
LB5ZoF0EAFF19IqF6vljmKli7u9otUFfvCQRyK/14zd6XwLmuyqN0FAjGB3EC2PJFrkicBEEP4Ez
KPEtShrzzIJIvBl2CNVAH8qcJ4X4tPcTJAUpKAfL1CsP9QrY74qhfcr2EUA3q9DyPkvTFpf9hqXy
0FCJQ8SJBczcrweA6sRt8MtVvxX7JHsT2qg3SSIDgcORMvDrPgAODflL4YgafB01cBh2r0YxiZvQ
NWOeR85dubMrdpW1eBSzeCVLAwtXnp2SgMvW4Y0iCq1X+S5DGoTjYskRWe5v5Og2/063aJjvMK+u
TG54tYE3FBsOBuNp9pl0f9mA5Mj0kPreIeEwMV5K/yzQL9nfzoEuYpflTXhw4l0XaxIlDEXkfN/0
zvV9R00vF2o+Zv20DDlnyK90S09aF5W8ESdvLzmSc0Iwbryxn4GTlAfyQXbqb7Q06hwpuP4QtugK
5S3mJ0heVBTz0e/d8J27QDMwmX2K3b26oQxYmupt5U6oYPVCy3EMLsOg7Hc1CnzG5VbK/z8/bRvA
KzIEy+XGOe3foiky61KlHmgiq5xfmnqu/jwwezzUCcust2iNgzFV0j8GE68krkUq/FWj9HAG7BIo
/b1cRfCHgm1F4dUxwAeEkEGFXUFVDEiWE8CjuHJBVNDK68hrEG+zRA0PyItsV/jV5PA3PABYZrOh
ePB/96Qi0Kw+gZU+w0sp46tytc8d1tB5l+Ervfl+JEvoXmS+h/nHDomfsnwgBuLP4poyi3PES6AJ
t3mwP242groUwiOr8iOuDYqujzR+O/b1utneEo4ir7FR/BVs6OiCoduV06jbyaRAWqxgZ4JfX7CX
k5ooCyuTjrSoYnrwJx3TsoXlQuBBNzlelHUgDgN7hSsrRCH3ZtfpaoyixBykI4Lft+nSkn4tCUXE
LImGgcBSUI+7Pn3lqa77Au7QUeWuVm1j3Grimlr7RReWnHH3cRFChxf+e9ssJdPcDMKzQD0qaIT2
euXlFQXLVoUcUUF4xnF/pOlI1GijZUrKFvV1XfDJPwcAB8U0vhtkwu30/JgiepXIXTdd/pWc7HUK
7sqvfMh6vqAcY0pmg8XeX4dJG/P4G87LjjZVmUHa5T/VtVO9V3wSpJ6nyr6sj7u5kOurUytb9f+j
vYVMLAqlAXHfc4jKZFnvZv5QG998kRP3rRoPlweTYVe/JERSqk4A/Q1nBn6gjT3w/fq0auVYhQnU
wuOBxciUALMDg+wZuilEDvX2a4dD1t+KfACAvYfw3inrQzhac07SfgbrnfFSF8oEZR/9IiKc3wWK
q2/pjocUoleGBVAvz0DFYuZ1CY9DPk+L2vmkkGy/eSL+PNAnRLpAawy0Xca/B2BPJunhHz+88Ms8
gumi7g773u+XSf7gKE0Y2iaQrBDsCuC4eArlwXUBGoXNCuTiZzdbZagqbmecw5W2FFo+hdFM0DSv
Tn+p/ykY4ezoMSy25/LvMmuvaHrjp5zzMKoF2ND/jzzGJGd4LZs/2S9poRgNiQ+2m47AXx9z0qLT
B1y+ZgdNHIz5x7Ah8dQDo/PfXVrc3gGUzvsAXQUyt/L2L6W+P196+ohvtjxVjcQgpaXCbZoPokK7
Sx9M2kAXC3Bgwnf8WIYSSqx1+/3aVcO440KXJi319RylsM/lPqUlkc5YgCIVVFo04j5nQXhQrhgj
v40h/VTZVVEaYgI63be4N37D/rVkke7WzGjk0jIAVTa6Bz3zFcPoLeemL26uO+05JtT8nmBGhYLm
6XX6SgidR2Zd5VNpAYLj+YAxZ2zHkzOLNbdSQOumR4dMH0g4xmkutYifL5CAjB7jYaimOTHwYGTL
7aBRRlotUKBomwQvYf768Rf2aJCY1yxAPSxBPSIcK2tcpkzxsoY8FWTMOruzFC8UzAFKqnWwttVM
IGH8xcNwUQu9SpZ5ku3lz24NiBZ7ZKsMgazAr8pv2BJhsDf5VmwxhDZmpZi/HApjcpkxFJW/+0fm
YL2/ztNzdSsjEsA8cZqX6vdkSv1xGH4BLj6wutXKQaSmBC0Ip3oGd2vuoHTfKnn8Wfcg3LTdJbsg
811nb0Zv2fHw9UEYxxIJGTkpCYBJGzSx/xNdlFNRZyvo9RPWivOhvnXsDfLMcckr7bzbuIFzkcGb
UZhQs9Cnrnz4MvFYsubSlhWfdZX2DBEgYOCpCyIEf0++8LaQAqqLe6pI2vMsqQO0+1uT3vxMeKSe
QH4pARBHLN0AicBmAuTqIPvRJii/Mf3vn0lx42VhdAiBlyE0ZTPKSrCgwl5fo7jgowsvT+/rXN9t
+SDkPE1EJKcue2Lo4YEt12piE5+Sl6ZmqMJ8ibDBD4xKgZGbicS1MmOe89+6Sp9CSLSGIr08Eq91
8jFGW3uMec2G3kVHN2rJSvrVmEpLOOEE4GPhm8nSgXyiowP3nD8xufdJ5p46g20iVfvXXdF6V3jr
ja5m4aTyCM7705eDlm8KX2CR/tKc654jtjR2nvFDLER5tAnXnSoZRteVrJ5mRlz8/Wm8I+C7XONq
7yF+zyJ9CsiBjdTUuyfpR+j+k2oZcn7bOrXzh/6KGoxmX1lWujLxotGcBnwJDORAUL/1qk3emuRD
E6EbNua9vo91cphA/rpB4UN6J6YymcXVoygqMmnZe3De9XenuMVdYGfY/buMo3ZxEIALnc04etPv
VQ6FmUILoMizJ3d9K0xOlrb0RGC7AX41RCqXFvjhYYedSOc0CdDiWe9r5YPAMYcxQKwqWGTU185D
rLLsqMtAYMlZShi96JnHbkIb6Xjpc2jMULKVut3ZWAc6BocoI8k5lecghipATRG8txNZFJ9IRBBa
JOQR137cGwpjITPcOZFtz7sbRCKhjgBKHJ5xjHZWNy/ToezgbNC1538zkFkWWMw7bjm6y+wtMMdJ
3Uvd10/lK+CMBZQGfGvgPxtbp3KDi5BvENV0FdpmG65gBTMCmA/G4K/DE3fHqyWqAFRvGsrmpkPw
vHQQpEe2ZFg81wEbC3gVqxH0/Ba/MhLQlUBZgLttzSuhSxTqjQMc0hazwxQMPYpodMDLyyG9OHYF
Cu1dBSQEmAfJXii2BD67cyL5FibKL3HyBHFKRUfhFdvqxqbm4GwOYBEXMbk7oyXesdW4QczD4FSQ
bRdGXVdN31lXDZ2210CHoeh2H/QjIDPCv4aOTPfyVhWnZdbl7z8zdZGVyH1Oh8DRjL1JCLDcHu/B
Is7697L8N1R8GcW6ljjkCfJA2rLJm7nuY6wG94WnPm69TOKk23H8ikO3IyI+6HDXLiICukMGm7qt
SyIcfygEonNT566Q5wrXl48184VyctAudrdGyVeE4jsBN+MhmxSZK5XljE87pUVBrSAxSYnEPZ4I
Yxk6KRCNLr0m146mvUJ9bUfLGpZ5YC6ST3eVKJpVMzt6+5/t+/rYE6ymGcMwBoZpkUX4JrA0e9fc
6C6W0g6npoCvH2LPhUhRpzwhZF3B36nUaSQVbg0NXRKTs3Zthi78WLvtGAUh6ekr/4SiXjTumVuo
Ald+iM52dknOyy2kEDSCZ3T12lJbyakWpMyF/J5rCEei1WvD3oYfLq37ojVs6ccD1m0DMDaGVHK7
6fqh4/9EozfOMD9IyrEzCMHspIOI6/VQZEcTYCRH2nplTmQXFRGMyIO4EnWjLe9q/lOad1MXXDW3
R44S6TP6vAO/IbscYsIFlmgNClpI6DZ+pwtgN9GX29RqQ8Zg8oXQ7Vr8cQzEbtnuTuNdXoYuny19
mtnTftYred/k3sNABx90xhkUGQ4lxk/1wM2E54PAb4vA+hx4u8kHgY+M0R/Xz08UmxIzH1IqznPa
n0rCOKrqsSqfj8QeEp1DyvoQQ4lJl5RoLRSV6OQZnNqNBXdsW9CNteYIAU30aC+OgM+xdmhV0Dzj
ft7BmsDi04oj04RfOgSwYWqTsTW764wfMXnQsi/E9c4O3KNljZlC+fC3plm3hFv4gOtQ6VCxCwlq
dgjpndIADlHehByCvH74S/oKbRcMUP506hwpe+Rb7p532brqaJY4jumBrl/2ayLEhIiNqCIhufCS
BoJG93rvYwUTOoNY8/2KuMOG1IAiUbB5zlDWmL7JRzfhPBS26reUyxD4BItQo2ivcci2ulBfR6ek
0LOjDzX+NxqRcRqQ6aURga4MMptyTD8d0xCUqFgA1Ri2j5gd6Dd+tvf1JYlDTtQHy8lHGEhuhDGV
iADABq/cmKj7qodfeaFF9vLnJZBLAMEXjS7wkbi0mtiK7/4mq/+IdaYnjjOYGr6Fnil9Z10MElHg
hADwHax8F0fy+NN9LWz0zvjlNm4B5jRGMUJiS2moMLlU9L91glLcFAxIC4jT+fR3dLFo8RmPL1Fs
XrJVe5FuLZlkTF4T/deOEiwMeDvRQDPIU5qQTWb1aJg0nUeXWnPkY2ZZDuX1vn6Urd9nawLNb1TY
7iwVDnV2Ifb30C3pTV5z5cGQzxiScERvrPVEX4X0tl6h2fUsP0Km4jEHbxWHIwuplwkXFtIbMV3Q
bAFAPytYTDT8b5aH2HQKSp71vICjj+AjGKYygiDzGsrbZAeuYmVD6CfNEs5B7m6iKW0N0Yj7gY7h
/lgf5Yv4MN/B1kvoVQNHqnWgh6DdTP3su18cQ3lWdd0cWiuDCXnoYHYSReZNPPS5mD9M7U2tnvGe
Kb9VuBaS3Y/NDbnrvl5ls8zZ+IKnWL/BFZh6dVphzfPs36do67ukAtTiS5Bq6tyLhMJ6uQPbN8pu
T0T8Dd2j2X6zoNsmR5I6Qb6CWlHeLZPgm2OKIKLLwpY/8FkYkxC7HSgVT77T5AT+YhgEzO+lYdF+
cGBfgaBPieIHKSdYhWPORjxozbnM3v5rNyopfQfgUwrtp4CJaN6CNDAWiBqmNnle64oJet72lWKr
UASqJqd6tA8NFHvQPNXL1jpx/3CGuwGBw3FvpuD9gV0SjUvjKJFNGGnn1LLv7Y/ejxkc3MDw/v60
3FogSnvBS98O5fM1I+ZUlJvXpGfus5QNWrxmt7F+7qhZXCRRGOmvK6pqxww5p9Zz56Cfl6SszFks
np8WTa8GRc5FNCuHuSMHGg1au7+peS0wnVgKs8bWQXUehmYUwFTV7G5l4sFvNFt3P8hZioK/QKzm
kOJuLa63SFZvhEeCNOiK9KlNEP8XyTqUqaHV+spdehBLbTq/bfjU9TYME21LCbqrwf0ObhU1PBZv
KS8cpJrmOA5avVB1EO+GWJ3b8UXpcQEAJWdgL5fXzxJ9xBQ8XKhImyFrKoxVIxUrH/qeEdm0fhnH
whu85nkdVpSpk6v7+tGDIhliIwhFLAxw6iHr7bS0gStxuBu/yD+4/tNgsx18JKb0APzILxnkrRI0
LsPV2r8nXk3aVPkj8P2ccpRe7RN3z5/t+JWE+rEpd9NNyvN3HxDhAD/M3KCJiUKmEOvPM3t86LXk
boiRFkOYhIOcXj2C4/OMAV0Ag61kn056Vj4qGpbno71yoG2r/CKHoncJ9WsgEziEuRB5aAijVtm5
OfB8AtJ1IFPUJv51cZRCMKjKocOopQ275soRAzaxMjxgoQlOVrw7P7qH69fhKXzxIYFxB/ewtYmT
LnAuWXZGrAFD7fd4NlkQfdGpJBnP+66+66H0DeRfLnGLKyZFJjv3xdrehHYUXTqgsyWgpHT5Qktv
GkGZXlC8lk6fPNDm1wucZYmBikvxnRaPIaL6qn6jb19sqKNHwVXWW4AySEDKCk/lnh2oxd3YhXte
sHA+t20Q1cB/S7W7L1oDtleWtvKIW2ig77ON+ARVoHQIlAQYmzmh2yjxbzRunaSaMKOJ05O88Bmb
85u1b85kk6MbEZGX+8lL3o/bHrKWMiToAm9EJxPuo/DiV2yeAEyYWGOWdNJewbG5SRGILI35vhqU
/C5y387CW3PUW9+wJSQ2mWPjMl/vWKWRw3niDpyWeYYKX2cS6twm9uBkduY2OugaxzQa8smiXyft
yxV7EKnOcYUw76w1bL7mJggZSL21R/w7eBNyWFhBWwQuwayMr4gQpcVATzeMBWeXl5gorDIe36R3
jK8/+lHP39Iu6G8J+cXXRArOfEzSOeu8UlNo3hmGUprkW/+a4/otS5I4hP+YXUTzEu4toYMLaU3A
8DlPLvkKvholZpikkkBBrPxS2S3nJ6RZ54wyqU3+FFCq/MPLwkrTmN8QuVdy+1vZ/q+4ooMdSKIz
7LXmvmyA0WSi83iOAqNLKich+79QDmvY1mjSBgcISqX9b1I/i+t9AdUvAMiBlDT+puVVgKUpI5ao
0eLXrPA5K3nIGOlEsp0KH2aAjgfeKTNolpEN6kqigxxeG2Cct13sM66MqWiCJwAajlF7+xJctbAj
HMuj7ln3kOoQvaZoIxmunj8DIjO0mEUIIOoudiiE6DlO13F6mPdwTCbLQsZrEo+NJ0avVVl7ARCk
4KHN6HdSCmmLTExlRDKekipvZWtTXbvnIORgVaOA1FC28fOuEWiGFLEyd5A4NYemabWzvHDEJuOZ
mcsTKb9TwImEKB8tjxlTsoClx8J5XRX/Uk2qlv4ViysbGF1q/hgfKihbFPB8etxpHpicl3C9FP7k
Typunm1YiE4bAlXOkMvdCcgyr9VqzF6lYO5tBAi+W5WALnxXl6qmyXdhxLQyDKvJKo0uGlNNEfkd
DS/P2WXPM7vN4qUW8tfYGAWC9kF22MEFSbnqzp1ZlIDk4vIPWOZ7XAR/qeMyX5gpzCF6/ex6+Lhc
sfLj3wLnHoP0Iuv4EoUh91X6gp8w42lCF1fji+dHwKnmqj4k+AikkiBLtlF3z4FTleP7CreiF/gK
GWi5Aqw9n0wkeQhV90/QKEn4QA7PA55rmvp9QtKzcnmZjZZbeF0mTNiRoYJjKdc9r57Lz+CeN4FU
Mt1t9qiYk+rm2hufaP4AEBStq96DA8GxSg2oN8JEiF5v149T5E/SmJrJG7ydGLmWaGWo/JcqLaJL
GrJDIpEYWc3jjPpmrygJyy5Eyo+4RGjoeBfBx08MFF2l0LeGpt3x1u2wADI7ai/pAQUQCLrKs5Ii
7scKFn9DBdIpoFYBIHa5jgO/Ltz5Ix+LZ6bD4TxXd09bJCrqwXuTHAWZLiuS3LO64Cc7xR6SV8NP
qcafomjQOT9wQNLaF83liimbA4toYV4f/5QL7JUl3DCkcweI2q0yO4cF5lK6E788/EJmUPgYAT44
vDxHHWlllpN9GS7fUlEcqBc0QgPulKG0/20pjCq7TDVUbOLqfFGxT6tyhllLSf3pUk8NjnOeDYyH
tphE4PXz4oPfdp1BrrphUJJJgHzeFyM2CNx3ZgGGcu4dXxC/d5LcWvk99lg4897pWST4HNZXg0SX
77w2Bmj/BD/FN27PM+bdwA0xQ4lC7jDj6fwrb1rRUtIobL7vXGoOIBDb/SNqGE2RcogXV9UTm3nC
s3qJvWTiPZf1+AdM5UBATEnQ123aRkYRbB7GaqveAunz7ZfEQTSFZefVxxhp8m+BZwTlxyXu8WVr
bAkwdy5nDScB5BCJYkhXi454MKXY5kRLBYHTz2tXXKF2Pnigv17EjADCg/Dk9+CbPAIeACUVSlQc
S/V8qi3vtII5iYE9erbdZjy59w8Wj+mcsXxRaPDiOBOKFUP1bz7tiIHU0xswzwdZPd9ZpnH5PPFM
m5Gv7wOLxaWfYOZX4eg7l+Wz+eQ1pNpdsY8P+g93u9dSOHjP6cCwbJWwUafm/dG//dA+vFasEO/P
aLR6qsvZrnt7uAXa7bOIhB4sOK7Ib6gCRFrC4ksGhy4EXucXhcn2DTn+hzF5gVGMtGDjQKwMVqoi
39Gi6KZhZismZPwYLKiaq/kmcnbocVEoE6jiFlX9iOgRQBVmzazHv5c6tgMWzHnzmH92FcA53SxS
4YVPGHfbrbYJVktY/h3CGOd3s2zecNrA0JkCEDcudJekO3rw9p9yURoGxQ/Y2lfA7DG4TAq/p0Ck
43GqQzH6iW4r0sVaYZovJNGfIASU/lH7yK/mvpqPAuAbvuVj2JJa6tpvXoN0K8juLdZuvEMTsvaP
1J7LIOzJLg2nRzAP20oYClUIf4X21TjQ8yPicGe9jwhk2hd6+80bHfkpk8I9MV6KMQI3SQ/oyKPe
+zppB+aq1Y8OAjWLYXq4k+qkigSMe63t6pIgPKfLfxRnak0PJ7Xnen/6/eWmpWFgfkzYWcbenHjh
uOK38WHbkAUXnpGveTaTEAkQva34idwJiP3ruxkegUMyFDxI+Ez3Tc2S8psycxsXenALo9DimM4e
ooTNHWKW34Pld5XKofHE7LYzkr2U4NtyYUlSw3XwRli3bqvkPqn5ZFLpQipgcw2IT6LSkD2bb37B
4feJSxvtyz/BjJkPctbmoungrOLMA3Oy2EfMOI/JiHuO+JF+nYBRzck5lZ+2Ep0EfHrpB4q/d52y
/y9iErHc3CFTbYdyzET/TKXthWcKYwEosJbIKo3J/wfF9uVwM84mjNyAAT0gN3SYwenQYDRT9HxD
DC0a6VV+W4XXZoQcuAnjv2fyJbGUzpqAT9GnAIxbNebctbLQQmC7ZLZsSfJruTbWfAOCU9Js7mfs
LiL05FWIedcyQskbsSbY2HhRxpcUFVZKGmNGvA/OG4r2wg4aRrnW+xCEoVc2jxnFjc4wADzz/W1C
HKpnM6/zOQ7t6E8FB+rCrPYVXsH53ZCdEjn6dMhhaZAKcWlCpWRIZjv0u0aCfbbp+W3g0Z7BFDy/
1hVCVQ3/V0YeKzqB6D5tD0sxZ0e2UetuFe6KfKvEGb2b4V35GwWOUg1nP8RDaUiaqh4AfTYx9bz9
i8Ma871rWlRTUS2xObxaDmmFWA9q35H3dJE2H3aMgipfFGoZdA7x0TQddZkreJNmjXu6F3n4jQxP
+IYT3CvX9KAQbA4HqUQTrsmO1MDhvzWVbcb2hVJwt3mY7Be6ruqK3jTOyumhDRIxSiP7Sbe2kQQX
mSdrOPVL10a/VfNHJOiK6s7sqVvIr6HcyclzmlRhLOuRFFB3ej2rMwh5YWg+frWG5qx/3Pa+Nn8I
Y7sm+zO80A31slSoipjrM0URfmljtrhgV6gla8UgkqmybIwkAhIFH0hFLY7QQQMxqT8AVCjMlHJ6
ctvfdlIazxIaMXD+O6teDkOPtj1lIfPvIN5b4btRjW+gK3OzfewSc0f3/a5M/wP+R8rRMRKjP6xU
P9lCgeKDH2ukt8Hy815gCPFq3ulN6kqI6MldZvmlXE97PvluXgPaUkwUN0JyOTFBe2vdT14q57f0
LJ6lGenjv78knsQEW63UaSjWJOOEv4/PLaOJTJH9fwdHy6iYqBfInGMI/eQ9GiXnwxRyNq/qmbiP
2GINi9d5KBTOl4voz8KHItvtfSUuUI/wATxUTOWGKzKoeP8PwTQdYhfSuSg3LpZujWXi0ybCXHko
8qYNnnR28cLIhzdSVlk6Sp2aDTct7miBdnsFe2x0QyaNTiJN9b7VgiRPKqshyAdHxkIBO9KSouhf
IvrzgmquXjlQ/BzoYN6gw+tmtW1dFlxp37tmfwuI+upIpc14DBlkhXalLQpLaWhhSqWxoF03lEH6
9eWpHW81/PazmaRIbNujFdsSPd3GkkskQhmq1lB+DtCcMTpH56ijlA7p1xtX8NzMo5ynuUDuygjo
ef57PKaCncvt9r/9lkXCBl/YsJDcG6kPg4iRO8qlX3xD6NGmyn4jIc/9+QRvb+xPbTUR5hohaL/h
He9yYNtg1TPNjhv1MaNK1NTDSU5M5K5WMkyQNf1rmrxSicwaTkzcIiVeRNcAOp62IL27TcM/tQh5
dXWKDE0fd1QAVqzKNcKKRHp2VlFVcf7wwCvU0Gh3/85RTCoZ5Kp3+1BY/VMpAfnu1QKD3Z/hRJ0M
bYYaxopJJYDgOhxnCjKBgwT0Uu4kwT6ynCrc881/eCWNT7zQtyzWrZEbk4qSbqOka5xL8f6UFaUH
ldnNVhX4xb20v4oOzYzCvOCNWjWI8Q/0dk2V9TtdmtjtTRzaaKkW/kC6JodynaRBhs5betTuPkrU
lqrVquFGgjAJcyut/zcyrcFsiZI4ehm7uOzvJ19sz8FfodM9TkAjTtJKu2aDhQY2tEMGkmh9HuhF
Z5kwLtAzOxuI7bTlOsx59Fkkvbxhj2Znp9GkNuURa36AVuHNLhb9J0p8FWC2Z/nIyujXAwX3q/iX
8dxiEy7dBajp0xGfLbBa8Wu3iLwzD8V76nJTP5m/sWwUg22WwHlPzyH8uAuMfu/nDiG3vwZX3tdI
xkSJDj/N2N0WTTBnAEhow1ZIfSPOrzmEu7d+fg9ocSuSuqzkCluLbQqtQKEAcgnOkijIKMX0NSE3
JoMIGrmr7xdmoci6ApG++k3ZlhAT04Zdg7vtJ6/zX6Leosh895duy7wpJNoawztddPCo4NQHT6nA
9GywWLZu/bJo/Ix7S7BqfdUHGRQsG32hD5QvI7fewfqyIQTjmXmqKpUOClYZ2YUMpGRCUcdMgb4t
j7uPMfyZkIFkWWYDYqWhUT6fFhI2P+d/3cmDZoG4jzVSie7kMSXbfUOovAgWRn+NkkZASKvlXGHr
hSKBpPQXbA/44PobmXX7ASFZ19o2PQtv8L5442COt57GBdqH+YuG/K7YazzYHs9pQazJEzLNF80a
xdrmlXeYJMIBI0Wv6WvWL036lx3PHmFmj13IEiBtQL1mQViM1yVwcy7QvSc9qf91MCcHpDdmfo4M
f/Lcf6HyjK4Qge6hF0cethc1pqu485Z/76zgkYYqWsqBBLtghagF789r09TVWyY+UwmJTOsEFOG2
JRmmyqRaxoZz3v6v2L0rkpK4Y4WHLSNC8olFWjw77IoVuOq115aW9RtxnbH33A+9hzp40exEWEyQ
DQ0hNVDWDfzztJgz2E7cfy3ZRHIXi9mdMrj08IIzmYkX28TSrxxP+5/YAXDb0hkekHvEsUphcW9x
/fhK8JDlN/Wl/P5J63+8z+5TzML8t53iuI9rlrDUNrnkMS7pSFaS2GqmVrt+egGGqMo8qHU4CvJc
o84qCNJVBfbf3daEgAr8543526Af3UkN44HQHziJbPMJcqEgTxWDLUGw5EAlakZgO6F3qmPiUxow
idR0zoSPaC9921jVIacdWspkQ/BWWcLWxRVt9VDtcCHKFvYK0ZDHSFZm+t4UhoseFWLa82l0FFYK
n0VpGtOh0/IKpwhoowOruxql7L5LnvbbmwW3CfQ+wIwf1cNFZHFISNWzTwMMeGSJkNk8JMs9qEwX
Kh8ktbFfZXETTX99Gd9YUxDYy2cyOWsW1DsNGoiZJYevIE79+uSOPLGM7UF3/kglI7l4S1rERa6H
PPn8dD/r51JAlzsBPQ1rHpm3gZ2Q3CxJGFsngrEvpX9sWTkaIyRJFv4iRg8rF+pjU+mcbs6MKrUM
r1hReMhM1ZYwUIKaDfCYDD7mQqvPsfZsCspR9fYerGt6etROWxWYCdOn0a9cByvtrCeMd1eO/0M6
KyPjuhXVmmhJZcKrWDmhHTRoOT1ysOTnqnYBnV2lsjup63GNGAEZbt/LqM7K8MWRKGzSottJtVYI
Y9dkcMrYVdPqmwAkvVjzVyV7sPzT34peZSZqPjLMaRiROIS+h/dI+w/3CC5eDlynPrpxgjEuViGH
udAL8heRGyP5MKLoWz4Z3FUrUjM4pKlTqc8mXk7LnWPWDz5Vt3MgAmyGibgKzjk2mCLoNWOkqytX
mZrLIwLSonzcSmFoFmyaKMfRb+vlZM0yDyvl1WcRDj7t/AxUY8Oiw/C6m7CC+omZ/vjVbd3ztn3V
6I942J6XWW6RS9UZsCg3zYEPmsKmhZcMm8i9vmn6LQHAytQOTNyA7CUuBYFMdJ1UAjItUTCFXfn8
AsFheFd2bIMTv0sn7r6TJr+AOpGj1HQSq1j4a3Gqed30MBzYhXNPe1eVR9iI/aOA8r8ozrZHtKO+
zv5nkpEqMYPdlSaro0T/BP5RrTUPjoicn6AfYwZ9yq8fgoQUxFcDnoKLNfP9m9lyU+r8DgEzN1qm
NshA4nB2bYQKT5rdcAyxN6sC10VaUr8r9zlPsMhjCBDAGG2w6JDg4UG6gyVg0/3AuA2e9T+kg40B
O5sqMaoGf1eJreoFkwwjxwyjz0sUeozvix13BYV+BuYucmML80hXFTo361W6xEODnglTJy+KOIfu
5kVqb6UQwsTD9AkKGku7qN9negAo3xcp2/AoF8p89PLZkce76ToXZ0O4+aB6akXEsrDS4pkpXGnd
OvoWuZ/msoRYmCEVy2sHDjePhxIbsfTr6Ia3nquFPqrijNiaMfA9Wun8gIrPxmmm5wNTKBVH5GIP
Azfj4XDj4ot7bEa+1w9zARfX1X0iRy95XtkjCgChVSHXE/SDDCZIXYqq3OdYR/HD0q8Vs//4pKqG
a61ORh8G7RW5iw+mUWHP82ieFYsrdAkSzr03mRSndK5QxzG9qiGDr3EcvR2BV/7He9KPh8yl0s3q
pBOe1P9/RXoMxIBa0tzzEBmoV5e1LFS3lnI5pZw8w67N/HAs7UGxg+v76cHyquH33p6nV4Ujy4Gt
A3uAQqBCeTzjXz0AKRD7zmN1cB7CwQQZ7pH0S4HehBOWnFEGdDH8yHApSj36HYAyKM/1WN5inDUJ
mMiHCdIiuO5fNLmeQRSb/RXB/zDeg98OQG5YEBGgJE/15TtQ7u/ZiAjVXk9cxV8wh8knrlZhlsuJ
MW9c6NlzTXi3IYTPUzkWHSQoB0Wg+Ls/CP4gGk+8E4CrXFisMYomBpWADUB83icLzQTgwL3DZ+Dw
jyzKLPX2XDYrVlYp8bNtyMYPQERNhTrAxwCvo1qdbC4hqjlYH0saCOHo+w1qd3no95zYjltrAWUn
I+zhQxIZ0faHyxIvcmGyonX0MkDmaVFchuI/zPMXGsvFDCO2BvMRCmI0K7ZxAsALEVWqozXTw4E8
zx5KdTPxBo5n3UVHhmKLpi3Gr1w10fQ3wZgDcPpggaQ/ihht+zEG/eR0LvgqxVJepl/YOTwxLaFN
QlWLUkcDE05Xh6ttbRr4d8tOACn6kYGHI/JaGeduu1Sxut5obwHurGmZf5jW2NO+njMvKX7btiug
+kr1+7wDbS0/h++GSsYjWxoIquNPLGh28IIYnk29tXjxfD1UvQ1XQCUle4deqWIZUfUPltn1U3Zp
585l5TvzVBQpMFTzjoUhGwOexJvuUv2/7ZZspdmAFfuYtTrJo9qxJMLMV22l1zYPBy8FiIUhtEeu
2MWlG1ePocebdgFDZcJeojeIVausqdqkKcIjSjsjic+/DFtU+4wFD4KDWKtl1PvLAxLoGdwOoGY/
jydSsHaxLNdYePAdmcP9uJWSXN7XoBssuqecc75kkHnG5ZdEP+eBEfv8oeCG0uSQFsBy+0YazG+1
fB5SslCVBLSuLwKVN6z4Sce/fSg5mVOcNl6tE47Vu64CjX0oW1DHO60R7Oh9x7qfiUR58iPhRWoW
hTfO6AzKlVBhz7tembbT5wAnlAWGxheFf45hoGtbi3aYcNB2obNwAl6NPmD0pyW/GWME2jNJ3+gL
LibacnXvOOw2VlxdwWxXyVzJPv1qi0qWUb/5qynL69Us3ImxdU59Xy1K7sK2WzxaJMwDHVFJ8ip7
RrZMQf2lh+1YTVlj/f7JjbbNpo66aJCdZZNQF6Ri44QePsZkvwv/91xo1N8Ao8PqpOXooQzt0Ik7
SoMJ/R5ADXCDj98UL55w2f/tSHcinkiPzjyGAYFwBDClvZrNKOPhOCN4FN9T+36sDC5OhSkM85Ae
1pmruMf04QN46EznL3UJFLMGFdUwrseg1cE6r0sMJ1SV7MSQsbTxwWokl4GghFz4avYkAUmpQGO+
O/s+8V8gz2LxdqJpN4qzvSk1cN0hbFLmd0VQwo/CHU5M7liBwmT0jtQabOiiCpkWgLO+stxUGrB+
7AZuxNbz/KHppZOSJT+n6gBO3J1Q+45Wvte6bj3fnEZBqRNkhTvAlU3zg4oU/+Z01iX5QTzbJ4vm
F46w3A7kTEyfRg9aL3sIyls2Csev5omWai3vR7CzQMdZBZVXPEjbvdWhhbjH0SFgxZhamcPi9Jyb
BGkVTyLicN/PMx9b3oeyXIFH7YShRtObSRn9gzGJgGrQCvHUhNm52e9AX3OtUHGFW/fP6ZL+8q9d
iiTdx5jA9d7w+SKyoJ1SZn6ZtKDlu//xuVztCmCT8/7ylPrY/zUo6MPwwBSSJvNM15hVzKDsI0kY
iDsaVDw6ToFHgGpENvRWpkx+6WE4qdHUA2jd5Jquv0/wYwmScPUbHE3oyP8wFwt0fQRMWMY9kQxU
d7z3XGkB3zo302Rg+zEmwecdeNRYx4ueYLUIUiVMmZBspezBiQDQCRr1iJrqD0hYeeiM2w2d8uBO
VOd9Sm/7upapmNVxAZ+fdsxFhJeBo0/yKPwrdP+KNgzsvpAWSRekXi+Li75IZPH1p5qkZG/HsY9o
UVwEslJLopH7QWdHAxSckXTnzsgDcCaeWjgvla1zJoHeadxzIBUYO4ubvkKhY5/cUpHFWQ/hsoJB
CvGjyww1BkvvpyWOOBLCJskmaGe+Z3dQ8s8LvnQTKM1NYkZ9i25Ep345MUJULky92sWC7G40ul+o
fwusV9Qc6EQi3zBGpNPwHdkJswHei6oS1JiT68VW81OWmBGST5f1WkeoeKZjsMNUZoNhe8W6D5IK
S/rsVR1lvx7lvrAw69hM5FamFrNpg1DZ9GB6XKolksaUAsZNLwR2naLl3suZg9vBdsVvUFdqKVYt
6f+mh2SaxLJTYsmLGh7Z67CqTDb3Ha1Nsjae8oSh9AMjv3sXuvYX4B0zbjl45MIbY6nqtO+Im4SD
taBfbtZHWR4wa+PAid+7xCYkDZ+iKQZix7+9tY6YKIz0KC2PojBRGsTI1rh9ZFyyFt/19Qkmykpr
GhLyI2EeFfJV6o4ftebLY9ZiTPu6vX+ViiLlDef8YpO1iEypLhogke8vo1WhdMErZ0ZCNLKSGRQj
X5PNINWKen/1uG3LCsw9TN0lzNQxY8evfW8a/tpxmBpE47AUdrWlA/TqRdUOopiKrQ21QBSXbB/E
zrxUQr+GSxgT3wGODXtFSnykjgRg/Pd4PdZZF3RzFJn/PBI9VUzNxK68I/rHJlb9NWCmdNnMckj2
c/gNY7GUkQUfduUpF/QhIWKfaovjTiKCW38GlXDg5353+Rln+AFjRNzOUIzf+0Uf4r7roOIUBC2G
411KUjtMkhBS7qKmVwx4zxsHblbSKX7PFJJwwR4J3DwktrjpNsxzXi7G1bsmALYhesRtYjKIoclv
qI6X/ZQRKavesPHtBgbRMEz9uy86T7G5nAqWb3kuDgP0+oE5hXdxUJOOasuOFRZBc+S/4QX6Ys+X
GX2OKi8Go5E9RcexVNRD5AOO83aY/e2itD6PxeJuZGNsHo7bn9/fWKkvLda9OnrwBYpLVgLhmD6m
bn1dDRbF8DEKyETYzHE2ECOYIHUutcKniCrXGmjADesh1DuxBAbhm0PWT/OqwneE0xBNnvTiQGgO
57P7TyoddIzt9KmTD7KEcyPCLpvCKX8d/wzBTj9Yta+8DLZ73tE+wQv4UM0UyqvKJ1g912WLj65G
UZDzSfbeYIeJtpj7IxW8L4/aeefSsGKpupIU0uG8911WNrk7+Z5Mnw/tELl7AGr9ec8flgWUXcRx
uzQjoMMc/on7VopO0bldcuJRXfrAhvlZoS3Oi2+b1lH8s0FhLPrKGtQttSqWPbmLXUlRV3CUqAUu
ZvGzsPXyRh2v+iZzbaWPnuE9Y67/pXiVqAP6gC8XBE/XbgOwiI62bsjm7NSIf6CNTHaARViYxJA7
F1ccEB8l5dTAoQZgZUpsN9UICNeZKeXk2VHFpLEQs3nsf46Wt6BZTbd1s0AqCYr8iceB7rZ2iHU+
me8KLqnjC1GZCCmB6mgPCoddpbcgKflv94/u7l33PNmtnXLodSgSt1BuDMv50x/0h2NoUvkoBZyC
JEWQn7HPgcE8avW+W6LNVUIyLz1C/NpbGTnq55/d3USnl8GIlGrGgSoF5+s5FLh1UtN1KVmGUQd1
iORtZK0/ClPCWEFy43zxwH4QGF/WTTGnnTo7k3qUgIGxAR8gHut12wi/w8xWMS4VBKFRsPkFLObs
UjKVgDwI7+X1e9T9PdSThkeUVPsJdEeLAzEWK79XhG2Jb4NqooLRGp/5xyTGIeC3vR/VeiuhDKqb
7v6twXZYU7Dy50jZo0Tw2NJbfyQpgf171p7yNJCz6ec9j3OlgPIflwZKzYn3XR0ZhEq5UR754DMk
Y1+o4hJa3R0KmX9+4L/ayYyQK1PZzt4MTXC4uVKoflrLPfzr68HjjI4yQQQCzT0RAbGppzuSOVFZ
mW24JLj2mhomAjMWvJJjxvyA7xHPaRXay2VmDzLW6RlyF2dkGrMzlz0mHC1ZvaU5N8ooTMYNOC3D
kZyvlS0u1YEpr4ZVY+su19hfcihX48kowk7y5toO7v96kjT5tPoQPt0prpSIox1Umskh+pT6NpHY
WZtgMNnBdSRtwRX0G9qo5PVdiCryerplltDeXTOgsQgjZCN3ZkvBau1cDR8gX/ChzvaOE5NLYR4P
Jqg3XyQq4KPRsnAe/nHX2ZOFAe15LH3Ul1M6uW7AxnUj98GqfMz/i9EavbkzS01dPtLQqve6DEO0
qQBt8wcKP/gcqQ7twJ7b0yiqySrqS2sqyix5Ir/ubuPRN54ygVdXKkd5HHdfllDlpwfaIWJKUS2o
0luZE0ROQNpxh0oqaCTEZnRs8O0byO1Uf74ETk58dWErb9VcHvSc+tiOHq1QjgLVDCYMAH8F3g4p
SJdT50GQ/9+AdQL1rkgUCDck9hDau+h3muvcpMGnh1i2ywkAsngZOy8OM+/XegeWet1LV7NlHWRR
BTuEhnZPOps97QYtJ5W+wPma/aKPAVTPCqv7bz8e0+dI7YZ27ytjDvXHej+fBz72qbVAAKItJFaJ
DYKI8R5SQxg2VRNik6YevHSU0f0TR25QUOoWTWYygqY2T+K+0eVSzW4On83k8Yd/S1zCx42HtgpR
CLmfbBhJcBoojkd4FUC+pkvuK74ICN4seCyfvr/WGRIzYezgkLBmBSF2HT2xzmI1SYUfLy0e5j9V
o5e89pP1Eho6gb52Mt5G3twkkdd4f0rTkcguAImnzf2hWvZjrWHiQWNrpD10xVyZW2poeKFVhjvO
LRxocFj6829FNysXkLKpU51NWwZ+vqj0+T2xN8aeyEd1vcqIH5IBWH0QUibB0vR5jjLmUhy/SSgN
XgP2nm1SPj9LyHjMHtf0Wg2o6LVL5jGPVjRZ0X9QgsCbpW/0LZIaCxSRmlvltVWLiWitaEBzsFvw
6S4emy9omrnkndPVGfAVq4MAv7FeoXrlDFiYcBNU/i8wLt4LnzJ3THAx8PFjRPq8VtaQ0LcMue1y
FvwYrA1wN15jMsSi57oGJCvNkFzFF+BCycoAHnQ2+GJY3XF7pU8UOX5EgB4PIhzfw1NyLbxNNb3V
L9xqrln7LTrBoFgcUQYSCuhP/jH1e4pOnvhg+KuS7ZtvbLH2hcgLGB8MAy5dRjWnN0wMNy2J55Ng
gcC2Hgw/Ge5XjcLKx0nDoTAERTYFdVdbWS+k7jW6j8yEmsSgryrlyu02QEN6Q2aJFVtgKvUOT+B1
jEv8Zx/DZ50LhvP858w8nuxlf03gEEAJm+8X8a5VvutHtS5CBW6FLHociHp+IHe3hBZjFRDoIWdt
ZneE9+Lu8iYB71wtL5EXT3WeTA98nUM1u4Kk3thF9clo0ln67Z4uGahAUMVL0mWjzXwjwNA54jIN
yqANyaK/1boXhJQAYXUe14Z0e6zNve5vFJA1AFMV055+d1YM2dMxQ7y3vJBO6x0bB6HqKDnGQCeR
DZtUF/VwD97gmqW2qm1sQD4mZ02y1Q15hbJey9JUSwlUNK4ywF6ANb/6sUY5bA0S/yUYcw6b1WtU
S+yPUja/x2Ms3mhP0lfB8kihyFL07G2FJtEBlEPOThnIC19MPTfy1LF3wccABQXjYJgBpph8v1sU
OKVX5qNuFpbGl5yVkfkWk+bHMNt23Td9/JXC6b8WvzzVmXIONNFLRfJJv6Lxj0bmchcoKySGxD14
LqB2g0eQhDMjJEM/yYzPKXVZDn55Oniqjwqw9A5mYUqLOU6ol68psY0p3TUD24AgfuPjdZ43kC44
ayY8ZdclKrxf8Jsk0UztkPBlVYRfy2NM4PYBbFq6hUi6V3V9Az2RgoYOGa7o//WCdiW61gAKDn1b
Qgg/dhVz0SRsPxzzvncLoDnoDFuOjVCKxmMFLI8NbX5wiOPpz61XUWIdVagv9Tiz4jSgx/mGEMzN
KbKbI72ngBY+1PKrMgLoyLsPMBDt1me/+oGh8GHkIWQzUxiWrRq6S6tUzwudXdC5HDcxLy0v//7f
NWEcV3vxFOslfqM6EmdrMiAEUf9TBXRqVWd/zx+Ltd/6TPquQNc49V5hi1TLVCA1Jgj23iLz/vY9
0idxxrBm2BTrrkY/ubiWWhO9Z9TNwfRjk/a4VYau1dEgLHxzt8UdjPzsN649SWI85ktqb6IV3/C8
Kozb4DRc1LBj32pUbMidFp9LpnbnvZ7ccP4/iZAbrVm4qXqmZmqgIR1asApFRmKJ1byIY63mL/tA
wkinDKiPvL/En6W2HlvTYrCFVZifOUDPFY7wVtYrHgk72q8PLx1ckAOV90KU5/cgqi7q8fJe3XYm
cITktjKbgIWPLs9+wqPfwAFdgbNPGWPW6zoLR5gqhQMlrf/dzDrZdcur/+EmDwS7u0m+RgljQQaZ
Ycds8OIP8PoAW+IB59m0EHUH11/pecNSYmgaTpJpTGDQ5wlkd2SFX3FRpAaTzTi7QWMMojS3huTP
lDhEgSXasczYjW+ezZrrCVvo7DBhkKeFJbNDcuS8LLundlXte0aG5ximXDNJQHnMo1dJCDls4eRP
9Ck2Wvkou7XHQ0SoX1hukpq5Qdal2UI+/U1D+sd22kIaMl7TqJmwGbphbJXQBFB5ACbNJBLa+nLn
kK15tYuyih73KAlosV5EW/AAZymLGzWLzvW74aiS+vvLdnBtTTJ5RbcZrRqCBggPnTieEOpLiCkS
t9BekTeKhUDjJOQmldvBMpuDDobokkD56YjNDLk5Lvn+1E2dXyYOVBiLbM+VkMMnzATovQw3ziIM
OxzgBWE3l/9sPNSiYKrut2UkTEJMxRkbtWQ/l3GfiA9al8oRbCs6zaIE1bJCMzCtDGccXRvo/DhL
2nKzIdxDTfNBng4HviuoaPURXompperO3Vh+j3I38j3EJBklpBqTQJmDZK0NbCK5TIj8PGYrVSUr
8Jdz/XvbCtVEiQBtj9lEDgB5zncZAz9dFS6GfFdwZkE/dPW5/l8fI2SEgRFdfC99wUBOH0y2bQ9+
MTXXR4+C4H7SST9g5ABT2cfYSljenUuwhhUyxma+mgVnt+rJ1utpFGFm8leKhF+Poq6MyOjYtiBi
iR9TLCAZDUTX34iE9PRwBUrWKGhoUJg/7/K8QGTCmfE6/UlhM4ALMSu8IT4eHMo+vz6Kik3F16sr
kN1LsDq2jCIZTkqqv8/TuXTE1bqL0KdSL1/CrChIt1g+bBHROIJ0A1AZZ0kkDseGFPodWJtefyN7
oKc6Ropn8+Y5Cvf1jXL3ybG8eRzlFmV4mb5YzvWULFexje6hWY5vGVRCyK1cYUjIk3ZUcZvEq9au
boGupVtjxQS0+vfUr8hsCzYV9aRjuglzHKdsrVQWTmh8cqo+IBFYIo4V22VNJei6y4BArYapvOmW
Oxb/g/brgR7MfMFeEzfAwIlhWlskbXVdzrn9g9Es2RE+1A4KRCKMfyRrfQZp5afgN9S5riQ2bYV9
/w2F9+ivZjsRZXIyCbtfpBtckp7LaW7qEPyNLNtczRgM3lUCrNT7eCT42PphdHWyC9lN3N+vedig
MVBTrxqxJMvDnDOGSk2GJmvjLvYxgTfEcZEPCGBpQQWhHdqfxMgdWfqvf2SV0mdX3XHePOuSRYUX
9rvvDTobtk+6snKZd6/Z57GZkRhvbUhWRieEvv6DnYbXdqXuRHvaF18pfbjG2LgV6cojTh9GrBpN
BDE/qKyY8AqiY5bh8JE7vTjFCmlADrZkbKY8QTQNOX85b2ZIe7m7sRYaqdrEX5a7ZkMoOHA+X4M+
iB1OKJXjHUTjV9IGOWiO2aatjM0mamdmS/c9ZzD8scqiHCPGpGhCs2Ah7UBDO/+ayIp7tilWulxz
F99b57aUW8VJCYIEf9BR6G1b83PcZEULKAdcfyrkEsgR62lMDNaBofVoHFJ+MmVOS+Hd+ssODU9K
JunKHnfj4LpcjYdOS6qiLDsCtG4sWpyAoCRNJKxdes+HkZRb27lt/qOo6ca7Th8I4mRpbPygt8+6
F1Uuy8kRl2azCP5MMK2TNMxcBtYHvrbmi0GR4AdFrzivFuS/N7FE2MrdnIJq8r+/q9fyhPtUwBq6
RXCgvDlfFYtFHcMqXN4zRu7ayquTSgZNDmTe4khHtAx6XVxHTtleohSjX1L/0GWa3/H2DwgVadDK
/MjTNy+weuHk5TASPSBWq9dTcGc296u3Mm8ChC6AJtg0dNdZQB9ydugeSz8yq1rE7qR8i+TCcNuH
EvAc6Sl3Dt7QsG+r8WmAl17BRH3aO6rHZzZOkGXKdKc8+AHDZ7IV98hU1Wx66w/DSgG5V8zF7Kbm
sOZgxRhtO4TXiuSoBx3CrU4rQ9v1kX8HBnOEpmDdv6QiubcwLMaUIBaus0uszgAnatE4ZWheRDb9
nSzdrqDGhKQ2E71eOj8ZxdAirPwQV8iRgDdxPC8atXNF9ihYKIDNXoZFVyBQqdNHUPVLpy3JEeG1
difjfN5jzHPXb09/u9DsjtvlqRYg5ADnD/KKSV9LS3Z8gXf55ZRuJdJdM3lFGIVblUoVZiv+F1Na
I5tjsbQuWOvkbA7slsbmBlsG6qKa37knMOLjN4RcNAcXZsxvKPZmHzItcRmqiOPWRvVetqP5WFCE
3tyU67jx4DILySTP3AlR54xUCIyNTbL89BfuqQb+D8gjPeDQNigXo9A18sMxiD4ARzBHVRa1p41Z
t+4Y3imOEirhng+fZq25tFTowFKuX1nOfThPbkXXRg8INHaYLMFgksjaFmuboNIWLNtfuBcVEu1E
3yf15Bt16KVQwdTROqaBQfii2S3NdGR0xFERDyb0DIE0AmV3eKRsCLmmuXqa026VtVsPJ4iiCvA8
pTlrBuAYYhpJ50KGAqfVjE/o4/uGRyW70VeBJeeC7wOhiKJKb1/85iV5HLuRozmmnh+ZWQ9JbDgC
oje9fualrYUFJ1ryudQLl3oPtQsGTHnBBmBnN0Lx6QjaGNpymcy+hy/+3YPOL0VWqusL4175D4EZ
+cyavFFePHQmpMlrITh+KWCbEIGXCTJrtrs7ihdVU1m5jt3u4mIpwUtAC3OF1BDBCRVNbDkQj34G
DoqYOM+TnWSQ+2c8M4a9QLxXkOu8WR7cgIxiOrsGJPd+b9nFzo1cZ6O6NyxVGokx36OnouM7V90O
XAe30nxQ+IrO2rdU4dfZuA8cqOjl+Htj1wlCUUpgjub07tLqbK4UYZTlb/Ley6DdBvND1MRhux9F
V+t4esy5oNF+bLnG+L/pJuYOWfXlziyNcglYpj7jJQw2jLnVFskfdb/dB1Bt7rGRVzh+38CrA/Bz
3fi03/JVl/y5sns3mz2LpncoS4nxPvBjoPO62quMDcgFKU5SFSrdwJruwm6BC89Vjc9AoYnnyoZH
DOCdzy6IVKTN0shHk6FTjdOiaaQBm/qL7/jz4Vm4+Daj9o3BebduSqZPQZoalwzMYGYgJCu2FmPJ
fZ6hNGVTXd15jZqrfhgAcHz2ybwV7P0wcK91/18JMm95brxry8TuSBX89lyIscsR/xHE6GEVcON8
zr/XEEaBOU+iRrGvzyDIDU+pBIqDuK7/81nsrUD5XGEZzPqF3zIp3ojwGsrknzvtHXSh8DXgj5SU
QVvV/mJW8DylKFLeiED4WALAVtJUvb8llgjZ6FDIu94sOGt1zdAggc8EzgVULVE0HVTStK5M/H32
kg2Jam9dxbFNV0OqwcEnN4dX03JnT8QV+yQU/euFBy5ral6gB6kVJnBk49Ugi3D9hA8iu022VpMy
9W4Yg15fAa0fAq1zcZqJHzBR5wTutX6my2NTR1bk2pHi6AP92Hj1sshjih7Rk5SAlAwBeGl0wFnN
j8XJK8wmVlj6Q46Ysd0abbQKAr19o7F9A9U4zqf09OzIyVi52yAsgfDdEvj0DTDRAaiyJG2EDm7G
OJdPsCPR6ebGpEAmEpqYwqikA/dQm8VACSVVben09rfZ5rwJKddpKn1vuQGQtfF2tC5rs76D09de
1mgZFHjCd63qVhhqFuKoNApsRQBEQlSXktZzTSg/a4aHb/E39c0sj+Bt5urhKtEjMx8tyVFZtoiE
ny8pRmuWWfXVlCDpp+g5gxetzuyS8NFRF2Wah787i1Kzmrh6UwihiWlbJyTtMmLgVGKp97C/Q2E7
LFWhbrjYmYBIJkFRn6BiGfTI1tEUvVx6OPOpi3kSXaooDvGJ7pX54fd4RIaxpNXxkoVtVL+HUCLW
Q+Rbxl6gmGSWam9MUADHhL8/p4aRGRXP1P4NnB3ihMZpYlwLXF8xXeBY1MV3xBel+wqbbx91OVC/
fo5mx9eoyUiwBSZNLmrzmp5Pj9fsLBi42JUqIvPMBgyFezCA3EkUwapWUx/9lHWY6DN6eN19GckD
3v21T/ERcBX1kysI5MIqLpQB2AlRMKW6mWpzFuvUwUZzRUE/X9/8kmfRaJWdGhEIyHuB4bYOQf3P
x5MA1AVUtJEoA68/HQm/kTc+PFWTXvlzmTFis2OrwuclYinTtJ2h12FCaFWoiTunw+AMDGyxrquZ
DW5yRx6SDDPGCDBzhi4FkP9fjDXZOxrF8XjrA7mWbm2xa+KJl5JmpsfHGoBeQLMx2fyCN3zvJ7N1
3Rtblu1jzsQGlYJ98rstRJL0hzMpzsv2XDPpR5ynC8cFkVuX2nFAh/3ATugD94+/U8S+E191rzah
KHc5rFgDN9JcEhp5vbrpbYF20e2K1hswnFVmgwOtsdxQGSPLTP1QjgydE2setVsFXSW24zXLzM9/
Td/6rrSRYA7R9j0LtVNM0QDspy2+U/XoXlDa4DKYiPwbNZ2mJY1nBcr2mxMWychTkuPWAkXlQCmj
jGIpttJGap13jZuDacdDKym2Y3JCo0dlCMVbYXGQGbh1E54jP3Yjecee4zH02mfrYgmDIn1/Ae09
qNuKF9CPZf9NTB0GHHgwnIDRiNwdWIpyAXEEPOpFGdDBeDjDi8u9w2TV78jMBBkganc5LU3XA/Zm
ZBPrZGp5SSFR7ev3d1twVzDs3pLY+QEBjcF2KkVLTiZbCO4Yfv0PptGxI5QnaNhPPt90WvYnoE17
uvQ78ZByd7R3xm8AgEx0c1ByN3feVhDTPWfpUzUQp9Q3p4v82TupEA6f2BAzEc/VLOb13ImoUzhd
5ZgdagQvFF8SRvwkAcZCtzsiUO/a9H8YG1T6HwnSfHD9cr0eTFWxpvcDZrnPMPojDJXr28uw1grk
dH3JIbFM33cZyMrdGxRpepoUSfWHXoC/iR/RvUdgTSzY5/anTFGettfgsnAv8qh0GGxtOjOltc+d
CNyuzzqGZ/6BATLqru4AJniD+gdhZctZmAf+Z921X7M/JPGSCtKDPiJwnhxadW0124WWiPKRx8kF
3sNwSRjdHKR0/IWjDN++3eRuMc9tPVeNgnY06av2xiK+oRUouBdueTYx2fj1S2jI/D+WxkbaaX6I
M6IekfTf0PBDV/0Mpr27HrdgEwyOTXm3BMlhf2bZzyK7DK5QxqTed2VGD3IGtra4sY+FQvmMCYYc
a22nAmQ7nHG0H5dFrAVcsqJ7oH4GDYrBSyJQ4yCKoO/4zemW0FbC22yAVVXw4fvcug1L9i2Iq/dw
g9tDohG+qLyvYd4YU5ZKjJbRhA+FIbTRa0Y8wlDITLsMIIw8PICj48xv/PMQHbO7QZ4U+M8Zx8gZ
mfUwTjE4N1plLrN/jkjehj86lYi0z+peeRJdojVCANW0WJQ5AP5rVEjKj4wMuFTHicvS4nMgYhKr
8dbxQk3mNIXdMNEQYmGvM+Eqy8NmLE8LqJUlGsTxBED8cEphmhZL99uixz6xK/NPltBddbiaVGc8
gwpVvKuwPU2jJ8jQfkTQzI7n7reVylCZ4GLkyxbJz93qRkA4lEay9bdL6UV5x3ebmUuF1AeRrAuh
lL6KEmoNMN1DnxEks80OwINBhGH26PKHpjMBxeWY1JJZSYlyD8tOBsj6M3nMykrv8nMDZFvpSaTo
THlOs5Jz0105oM8LUe1hVy2f6Us5J0sClM3O59lqFSTkg0TPZWbrOKEyUOObbOtVsoPVgocRxGRM
euRYqdCWno1ZIV9/NYmRWOQd6BWtBa9R+zl7tljc+leZj7gwcpfQE6SRKAHoSDnO8+9MMpwkBELD
+QLqysWhSJp2bBhJn91dENZLNehCl3J1h9BNQx/9jLdXrEzSCM8oV4Zv2e7Dc+i9nz5VF18+ciia
/n/4jR50XkKwMYknHWiZRXiFCllY09DMm76ZAk8iQynTsYT0XHdH4SkdEAJZjtT2XbRbcfcR8MkZ
m/JNnHism9M4B3xGVhQI+AToQUQN41YGVtbyt/UPPAL/M8Wh7wnp5DOCcf+yGdGXGWUhJqO1LNqz
iKeSoZ+mm5pTVuN4RFhbtnG180au8oy3adQ8OcqnzWgIw5BEbzdUYB/CWGceEpEqNtBDiH7U1PiF
Rh1ZgIYMpVjvWTj7ydZQuScLWoB7q50SSpSAzcY20oCKhbmCqKy6XaSsQsGz7LICozY54uSSjPhN
2U5sVKQeTuzkV51j3rS7P6yN1t+ogKkb5t8VtbpSJpbgF/MqwyVVCS7Z1eFXoKoJPRmo4Vjnhr8O
anYR/NiMw+WegEAGJRQ4gyVom0aott9TAN4Gvhdf0zdKC5s9GkImDY05vBY0YPGdwqVns/VNZMoU
A+Xf4E2EPm8gQfs+F3PPvAbnw8Ap/uvGtbsZ+eAgl77mMtY+hbqGURQFYEPmxwYO3H1/LTXR/B3W
luoDxCD2DESU5Bgar1pDaDrx0MJpPyQDaL6ke6BMGdfdOSkvXcHagvCq0DS1WUmMSttyiAM7cmbL
/789uGDUmrApiIHA4IGQ83/rfrGHxyJ1wMgEQzpq5aDRtZRshXJwhX2r8sKZ3eRsb8Cdg5Q0ZgIr
YrZ4sFGVkcS3AlWQEIJwUpD8GMBKEriN15AhD5afgiPhmn/Ys/ExqLmAslNUOWV7klHZVPh2SiMl
mbmBYeln1TmJUvvoU9hioOI/1nyxGmdsNxXaRxTgCmw2O3MfUzRg1n5xtfoNtaVSOBBRkdo6B7Nn
eztlSIkK406tRPfew4S6kq5rjeM0FuoWF8wsinmhIEHtaO/iPUK5L+7IXpBZMOGR2CXRpUmdHBJt
yvDQgmchrM1iq0yaG6I/dnR+NnMJNG5oQfCUgywRp6WNHsWM+DanH/WltEx8sAqL2ILh+ARVhwUv
t1U2X5l67ls5no+L2l3P3GJAy3k1GWUMlAEYf5ta+CL6jkV4ZsY/oJA7fT+LDM1zKoSOw2fj5IKI
GguyDfEJ+D7MsNbMVv/U0bhTmCzYBJUwzrFobtpbq/exA6uW8nUw8Ghf4/cyXDoIqJe8nwCCBLN7
sP//ABjXHV41rolQl9ZWjZ6g7k8NcvVVe6HbWtrucZLGlcO4wF5UiAfi3nW2yIN89cmrzYvcdJNL
dBDqdsZTktc0/FwS8lu/v90KfnGbRj18Q84qsmfkKTni0DMFL/SoMbP/zSlHL90KL3CKWepkduBP
2tLkKEki8UgjmAoQvrrbF9FfwQxx/doX5yq6cNy23ktPRFdtEA5yZGNVIg12IXHlzUvPBdiGWx9a
SbXXjCmfp7yIvBBL1SQIl48SAv7+g4DEXxWtMEITfwwOfXxACV4+sEf5vI5tf8nh3AtC23Qdvn1F
8z4vI+iYMA1cytL9q6K7X5UCM8kNEU0ZGTX/3PLQu1s1phvCvgjPWGhkli/IsOE1mv1qCt4hnnG7
ZX8fVgFSB/p7m53Etu3UpIfTTPI5XZg1zeidJRSmWo4K3vju6VugrudvsOxmjxpJWYfpoHrfuCVq
MWYWNCSVdJfKrBwgKhjnQJFT8iyWEfdrizK7aMX0zs5RD/YO2L69HpP48CfMrWZNsTmUpipLxN65
3zn75phBM0Ue8LPdy7Q9Q5VfIyjnwe0z05crV8UyTFSY/fgv3fnsf8Hi5T8aFRo3luhO7o/DW6rY
7hq+rL9eUnQt4scrYeUt0ZCvCbVpRhyqjeIUEW+eBxuvsM07kBfIhplXfXhxKyKUFiem9q+n7PuH
qChABUb2Pmq7nTqyfkCl8AMnnDDC0kE2GeLgYBsjaOWX1hMepbNunRretIgrSvctFN6fB0xKhFar
KbZiwozWGBF717awxhVEL5aU675l5b6Cf3pzenUPtTuRU9acyb27BF5KoYVbjQJxaXVa3+J3svFU
TkotrejLUaNTub/+U68onNE8BK1IgYbU9u3y+dJi6MQdipGjiMZw2ISpHGSiy5NQQ/W8oBF5jqJ4
gEneARbYOo83xDLg9Gs3Ar9SSKYKL6QjuIORFwStt9xRY0Db5HnzEmbGmcOm6Lq+P5AQMyHUZM8D
nVSL/lJzZDyM8c11sw3pvmNvA/yujV4Uf/VeZqdBxkiNc4CtCozWKhTEWy+Ptyg6jzsoehLZAnyy
IBZ+/oRyNpYjXio2mmMd/N31mK6r64aU0qF31+lsALbyMe7dbyEFI7ovFlhXiDQdDaNxAADEn9XQ
HOUO92kWI25wTzsXTByzFdcb9Za4lSeyBj67AYa/plQXAW8spmRZUwnRrhd3WTCMQXI2vxJpX6Kp
JHslHtI2gNMrx9ZQgLwfDBIxuEWu8k4sZ9ysQRxFa+vQgBfb9aOLRIi415KCW3VmsTjHzmL++GNP
lM5rok8DcpJ7Kn+mQri0i88QQ5AXN4qlkvEtC6SZvohElgv/wMA6tJ0JpJiD9mNPnuE9v8KUAVDt
hI6jNYoFLsv9jXGBLiss+egYhNi6TxikxvEDQimZX4UOXJGRbdwu39bMTjYB8Um0PF0Zz3zQ6dT7
zSGOjrvC7ufZUJohNCmEEBHXHQ7vFBpJ/1qN7R4xl70LuEWbOsd57tuqNwRALTwtZOtvyfmLsm5G
TY8BFNfz2xXWl1/vi1P7rnOP1wh+THp+CMiukxAIi4/EBSvRAraMOKmo/C18lbp+hGUsJIdoM6Db
Prr9el/djqWdEm4okqzC61HEMkbXtuh9vFGN8QVTmmiAS5tHTmsYaIkhRtjoKH6z6adPlD9olyrV
LXxBksJjDZ6Z80t6w6VQt09GkZq6U++FhXPRzH4j7+wPfmQ5MCXT/A4152kX75uEcUuL3Z+TFowU
HVQInwy+cfMJ4gDKgATNmcOKYiWIvAMdI1RJW+iCzYSkw1FMKw6RjkNup2A0aYx0WDivMOVW6g9i
pU/IVxxy/R4MlNTxK+RnSVMyQ6mCoRuuLDTt1HsTtpWwXLIKWHoC55GGFct1qzxJ31uyrEFJvinb
4SSx7hfx/KstJ270/cI4SlCwiK8m/t4c+/IA2OCoFtEz805AFqzPCHhaa/SvZ+WaxImXE+7mZyoA
ZXfzC7o2zxmoGulW5P/34NzNxpS2C5/g5qtM+9flPWhQx4Z0Tsjj+BF/ABZzYVdjCh5s3Qu1Bibj
dxLbgtkCcMT+YNxbXWporS7OBwXiljTwm23c1FkstTGGpxvrMkJkm00BBwUY29z5cYUhypS3lH/o
apR6TYhnYIPnyayIXfWD4Avb3NhxZ/9AKdRXrwGdte701EdyYXb/DW0xw0KeCQcRYkb9GrkLg9e7
/qcZ3ObmP4rA9aBimWFLkhhdDLaVTd9bhp97+csklha+Y0nEb0xZySCiDXSWbbQj69NwN4Oexy+L
q2woh2s5SvY0u4g/6E+89ik3QusfqQamvX88dMqmv1JqsnDA1oavnzlkuGPHk07rzH2ZZ3N6xfe+
kZq3inGAX0O4fU8YTWbXos1oUQ3mf0SVyEHVB+eQYeTO5vRUl1QvSDtCK2m1js2TKWeTyy2GO9VF
7TRFSgxAb/D/FxQxy2PvaifF/ujyZpDdmrhTOnSR+giwJ+IbwkUZwgixnd9Yjl/Dr8/h2tOC/od0
nZuhpt7u4eEAriETbImiTvgC4H2fpYwYivYrPo0ErbegcA2YOBNbjjLNuFMScNggAmQylhhDcQQI
HcbN3c3/s3K7+TDFDAZxEpXnC3WDrws2te6C8pPRkY8SYI8bMZwlqVwrAMwNyvzoR/JnHNjL6eD4
BNFNlHoo9p20Acom1aIFh7mMgZhuACt0pclIeJC7nbS4OV3ShNv1TOcRv5UlsfWNe44dqXv5ionM
2gFRiBzZTLTWqdZXNWkYEtFvB5kC7K374q4c7tktzOvRZrcKyDt29vN310snG81cqM0cAIwECgD+
iCuywdPMBb1SiTZjeRy/NqgVCM3tChl3JGLQqX+Q2sjEmoUw67+O/F/a9VBy4f3pifNI7pNpDND/
OatblJwVmyBrDxcFdTHgvHodG839xvHzdrAK6FmPyUtKSw4gjaije29VfmG0ZWBYE9R1zzw7FDjv
tSAZMjDztHV4xhbNNc8OHsVPTkIrECey947rB/oN4MgkdDfXvc+hvxo9/xxqfFKOru/TPW4tDvA8
1vaFHExoyXs74MnWv3YyRFSsaboM6Lbitu2v4OHpob81cyTob6GEGYa4v7BF3Of6oygPg2AuxnRK
sYfLofAVkjvrVvlbe1dWp1HMdOUlvcKeR/zMpj5NMmO9REK2GrmTjq9KEzHxj5i/2/AiyAlW2ej+
jWv+Ln0mBxN5Jv+EUbR9XFsLzRa0bqXBbFVsfppEOHwe9jOzUaYpYrATjPPcLucgQTzYAdNQBtIV
q8dQQ/YVDCIFb7L8ZgjcOdfiVyHCMq2MR8YMoPCiBwuooOTbQqFMrxRggbRvzQD65c/128Na+ker
dIMkHZ/B0Z4lwA6TwUc77FbgUIvdmPhRH8jColG5229zl/OjX5op/74+8Vz4qVdbfHZZz14QfIS5
5rMDNJ9Axq/R11A3157lNOWC+7GpaX74ynbfKJHZNXJNJhc6RdLrAICQbf+rg+gAT6+5iQKE1ZMY
s5+EcbptAnA/c1nBr1xn7hTO3OPRIlGCwn1fO9RfHBYCyXZlTKp7DSRLCyhN6iI0gPaBpr9Vti73
wEM7t8DEwLFOnPP0/exX2esNbbfVe3jkgcEFKIoBxmZ3XltCPB4kedaxPMeE96RVYNuzq8c0vdu3
d3LVGyT0LnxNN+QmoCCSn6Q767Elf5v8AnM5+rsImjBW3R2rUEkuFVl/tP5EbFjHTud5uAlmf2mg
ihIRpxKfhAuF3xATBEu1GFgLyMg9ol65ZAcxbqjGKPpssA8nx0dNAqEQYbmrgtj1aQvKOUAm0Axx
YSUlgi/6kFe5aQsR8fdd0q6PY/vSH2Z7jbQ8Be9WqPzyPLigmhlB9CNVSkfiUbotHTSlmXn9UZZs
xiJrhfjm4BBbCzxSSR4y+e/LjkiNELTJRFa0nefYerZiYYZrdrbrIf+pFGDRaPTuLGjsD1heVD6W
b0n4gikJuh9dN6zWD4BS6rogWI+Gz152LqpaSqTTmnT/mcBPTGgzZEWa48ZpBy5nGE0QM9b3gOzG
Cv72UFjxmn7HsP+vv7p5zq6EGwTH4iy/yByWBQiR+Q+BDruYhY7l3BeVgjoSu97+1dqLFPfAFXDP
wLgQs2EY4MqXA+/Dxy3ZJRVTpwjrzbRJW+HI+7bz9WLOsVG1GLHK9mkKk2odEmlqnxY2t5pdPwVK
lUS1leyx5qi3akeCy2iPbiM/0yMFWZD1W4AL3KBhNekUNSvkF4b8YYMZ/q7Mx76lXNbV9qJNRrj3
w2g8fwZMs4hvQbk2OJxvlQ+fGHNN90dR/caInlbPpgCH3afb/EsovOrAzI3Mnc+eVwQ7acqAOKWh
3U1AA4RGtD/q8vmzRIp7lpZeNAvNksDB8d3a23viZUVpWRfF2QS6svS7e2pIA1XcMWCB36CU5PnQ
QNYsR9H0GdPMb4K1O+ko0kOQj2wkpcIi4ePWuvcRSgrSZL1h8QajkNgDHddLnpW0SFwpKopiKH2z
SIQlzswqxkStloFq/d+l5sVXM6j75WzXn+q1+jiPU15CnY+yP8dJ0qgeNqyICPY3k6vEAFVI+njr
dY0vvPK8QLA6+FDVXZExH8Znxu7KlTdk1I+SburLkrpVDRSij5SSEz+2F0gfJRg5Qk9K3c+p6lM9
cR0WlqE/FaSdduKC+NkbZKhCcuZzqrvCYNWXdQIBglf4PvcfgvWk4BQDmJgWfseBctVxn35igBOk
9GH2EDBwrHHVAfgrC+2JgpkNimyqBOIGEcQo2tFKNC/7mGx5hnsywUh+LhfHOrujRPYifEAxr+bX
30M47kF3/8wzju1EFShgrzQmdYGkIsNqTumwfVtAzHZ3oQelkkzZBK5TYHPngpq2ShZCPER6iodD
RLvSfCv5ColTJ0Sm
`protect end_protected
