-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
JDUAieB2rFncIYCJO3fIFZu6gEU1OM2bBkcUoiHJuL+feuuauRWGAMgeU6n8bS42aAUaOUwEyVrv
euzpgZJ0F0dP6cNqDud7DQNyyFn+uFIxFH/l0TDkdGRX3G307/lM3B+bmHRDJvaWtWZyP/vbrcOc
GpGtvk4UXwnBzo+JG42pbllEcpYSfFWICMs6vmA50KqysybEVo5zu1ivM/3A/G+jXsX/6z8ImFMp
0C8FvxNJIJT1CGTO67vif2cRb7DW9FIDLADPqlZDAfnUuGqif19nLPGKnsP6+NeYNJD7SPIrUCh5
GdgyOozhH/Q3mwGpO4dVkEuq34KgFJ7CjIO9dQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1056)
`protect data_block
nz166GKaJvcIwIb/H5CTN6NrDmIwIQrLPxYLbw0hY8JoExpOJcECr56kOqBtdH0RFBAx7sNj9pXy
gOFLHnGBuE5HlHTx2l2mggHAC2Fy1RXDehfsFiV8WitFR29Ib9/528tbXIKdiJBCB1fTSnic6I0j
SdMAKHS57kYr4Rt39JZ6E/QEMjw7IGihFfrOVqbUgpgnYdjqFfTpUwsFK0MDpymLUdniIl6vq3kP
2q1OnQpLdh7UiVc+lLzwKxhrA73vxwuFD3I4bTEN0hDxCT3La4T9Rg/v/AWIGhru8Ldr1N833V8T
5tmwsoYOqUp6+keL4Aq+WELCx1d+2NGe+758pDPPIrbdLxd/FOcP0t0ra17y3wskiRCEt21s9jLQ
t8vy7KAeMmJkdw1oLP7XMNEwjwTCf9DxdKEVijA8wGetFSbi3vK8duuETQgj9SPY+VWrW4rF5v6Z
5g0hn4GIei81VIloi2IM6jSBiPeJp3rIbkhbRPVKMDjbrqlNIpnofxJdtKSCoqHNqyDnT7bPqMLO
8x9VxuLMYoo/V4AZQ/xCY94cc0U3iNudbOjCTo6N+BevTQBsMkP1mHDkm+IUe/Ixr0268a3p2WcZ
N/VXN4lWA9CqZJ3j2juIE4PEuhimmlOUOOlxIvQX+R6Q3Mikq7xjwHJPlDO+yDS7q8J3Tf8We57C
lZEYsv206KwO0EQgpEJbTghwlbEs6JhKm1cVF+94HZ4x/DFZ7Dwj5xCZlLPtGj89wAus/M2pjbcT
yCBduIJlCACiMsbtAteOBqV7SNGBsVKdH0vblgTNXPiZ29XJWKGFOFdzBMqA1NgSxvU6yHhrzVZ1
dgeLR47P4YNTgKyGVBuGd4TTEXJsTPx1AIICbD4ujg/ZvUFjROB9pCJBdvlxHBV57SK7VpUWpnru
wSZ+5baqOg+sOLLsk9dPjJH3FjfK00tMHiWQPv1ZjCYwXggFnpMvTT5mhTYhcRGhopu1UuRDEGxB
Aa9daGVQLxWZq9qLrdMk41qstElDbRVppwK+DlSDU24IDlnc8fjfJZ1BqJ031i2Fam8BcOJE3EHH
tqjL8eTXOaokjpft00UoCS/1i7VF6pl6Hv/y3q80Esf0BOOyINihmfuVxUE15a3ZJOMgXz6qeiQr
i/b6YdG4LVgt8JTLBlg6NRYpPvmdENa5IlkwZX9f2N3YzQSiokHA77T9bXweHujaYyOz/Dki7IP0
x0wiQsrN+UeB6//yu0CAud+iQvjBgep2d4pai2ePteqrSBil4jxp4aweadMOLdTJDoluTIgZm+tN
Hs4n/W8WCgR9bTnChac+WrTB0yuzYJD+ySq8/sVoEoOj1ZD06WZGR1ZymO8iGI/CS9Ar+sQ9vfK+
anMrERT5bMtbO0WEbBDneaqxEun80oPZRQ7LPAvA
`protect end_protected
