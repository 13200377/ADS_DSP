-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
IZ4d1cgsVhpKkhDJFzYV2mkpTgDhgZsp9bNDYevPbkSDVXT82PfJbhgiCeS51E2Vx5P3mXAtGAHO
FE4ZDDCFbzgGEQel+zoJrV6bVoQmPrSb+tJCvJ4JHbUwQKyol12zBWi1WhcYNmE0R2XHWP1B1XBD
nWKoVbJH0K51QvZv7ZJhC4pvCrozMnoatZsOJPyqUE0qDVp0jxMLqEwuZm5B5N1xT4HnJOoZD8AM
KXpubdfIXMVLzdns8/njfrGGIapp6PZlynp1p9phG5SGHTF56TrbH5ufVNCgOhEJ1fmvZFqRtCa0
3yriE8vL9DXnSuWN44YrrmmM2S85v8yKhPkPaw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10336)
`protect data_block
o/8sbXAM7zHs8SUSBzsL0PLlrU+CI2tNoN1teJgN5987Dotkyoiw+JUZd8Gf+rARNml6Jc8lH58m
osOK2v++0n1AgF471FrRQCE1Dx1TlIV0CuBabB2/zcWY3Mga7Gb3uirUX8wcqyNCxVlk0VaH/7dr
GKLUeoA+hKVDEj5WGUCpi90SXiFTb7f/gMrPeutLgzn98d3u8EW7DCOpQ3c3c+ErV3OwhN+9V0zm
AMkK+mJ6O8Yo4f2RMb4ob+WSw3Q3za5Sa8nXNbs4sSBr5izLDCSyKnigyyAOkZP1VnVF1+BWLfJV
WQbfXrQIV8as9/Alf+IAzB5bTcYPtqasHPi7WAOVOh0Tx8f7Qxvk/2mS+/ERIBOLA5Tc/P2vYFXu
CHZ99Z7owVvIoBP3DH6CV7JpIBXX9Y1YRFJ3Cjp9k/zml4HaPKmXa/oIvR7qmaqm+n5YAH+Oe3fN
RKe00ZJkaw+DjXbb+OOrDZbdQcT8d7BAPtl645jmQ8IcTcMvU/K4fMzK7SK9zwtqrcHkyKf7p1iw
IjVq5ohYaweKKCuoONus5mbIhqOKQjEZCElwgfS2s1+8TP7agkBtg0xyNauBKGm/Pn7g72K0iogC
JBFyzkwzGjK+mxChE/Y2XneyvDhmQ/GeAPdx54v+Zp/7JGgY7VNBDIquSIqxJ3YfpRMIEwKOOfFk
a0ogMwrqtA6hLHtuv6Wl6ssP3MeUjqhUOhBMvWCplUVKkbJv8zdTbJx0nM8YzGKsoD1EaI2dhDZ+
EoP0S9sNdz2g/WGx3BQorUNCdqD+PLzpU4hcsrY3KKukudKfpJzZWs17vEFBlZGfxV2KUR4EjV7X
MEeSNMRmVij1FWACmrRbakf9I7GETNcfmxLJ1k4+L7rzZPbcOfnH8ko+VyYci2JE9OlcmK6ymvX1
+9hLhyNIAFfn+AUmRDg8wf1esYgk85u4WXLVmIZhXOs9EUYIMNHIDp4TLP4/rz3mDf0Ck4s00W8Y
iEVDtngCKUDqiI/3PwsIBgTqFiHy4R/LApK945AJkjWtwy1iUjogZuy8OtaU3kyftVyFIA/9b0GY
Kz0CRmMoYLnOrGnzwQkXNylqgqQZD8rAdcjHuelirlXObl+TK+qVrKQ2Gc0dctTUp9yR8o9+jews
lpoeGvsK22cIqt/t9z0cVqGsI9niHv3F41w/V/gLLWTEB/uh2tbyEmWOm6oSzCcT2QcWrVPW2Ny8
Oj7203Vqs7u2JCqYfyGF3nHvugdlC3FW2hXJoM3pfvQMDumBTiJWcxe13HC5J68xKmMr5OLb5nEU
GSbYn/TjmhloFIe39+zo8HjrScEZr0Fh1lPUXwbkYjWxBiwrqsLp6K5jS1H2aY/6J0jsyJSmXiC9
RHJledIkYOs3uKWYqrOlvC+5aYRKZL5IUYuGoo6/lWahwloD5DtlTi35mRd7QnT0DHgKqbV25fKA
wRW3y+ffPbPtf3GnAMPL7ZNmnZhqaCoaX4gDgCtSgk+FcMoNUj8+6pMb4oZqPBlKMLhlJ4N9FYNq
pbawOKmKoAKTJIHSfb9/3d1O+qZvJ4/gyOTNpYFkdXihkneFu49ij/wJAoYyU2o0uM+480Lu7A2S
MVm/PDHcGMhusbGObY1lKvsTFhaMNhIz8P+k3H/wP7tzX4wPOM5mz+Ah6Q5Yfu6Jiy6tgjD8voIC
2ud/xeQRnwL+mNp7T+C6iyRycKbjoK4aVQLYaJJm9qvQDQ9GumLj4X1zsqzW6gPMEYbjpUunXax+
ayos/LgMsoOqJafPGhJQ+VLibcgmnKFs6tBxOfIxbQ+qwVNvGuuMHCMNPT45OHlPZyf4u5DTIZdE
6oCiI3JeeYAto8HfLyQmhb/Uax0gURql8EdCLTbd9PzbxugmwHve2h5QVu4QUxKZS//f748Bg+mF
8cP/dODnWEP+QURfTZ9VioskN30iE8YouKL9jIp5mvjBspm8GKxtu87SrNAHIXwFs3CKI+8/wqk8
kKzdSJn6D+8PCoUg742FBqK6YuJgFqVeY3clSHre717eUwfZT090cn/Ix25hlF3q1hTnzN6mxzkm
+pBgh/DL4VauvX0Ts7N9Xr5HXthNs2cPgmC71DboBrSb0xFC+XBjq9KHabGKaPDc12X3eLG1+W7S
abTPlhMO0nYRDVNf7f9A/uS2bX8H3CjBVpYBHu2DEksHntQZ/lXeVshm0649XqvRuMSXQk/xKPP1
4CYkJkSRGLOOp4Maq0SP8cG9yrv10COujYVtxW90oBclauSURiCHJJ7VEfNCqZVYNfNfTGlHMX0e
LOr06OEjGqK/OWGckRI+GRdoySbGkrzAxnD8v7x1JbvhwX7m3/sYx5zqGKGA96K55mDsjO/cJyW9
+5FcdEhVU0sFzNzyreyd2Uz/1QiFCW7X4euxH9u9dDUC5Hw+oab2KYVlgXrCGkkik6L5xhzr+36w
ouwHvEpWxh0OwHmWN3LWOprelA3vDLqIOIEbxI8LqaXBtMJVqYTqB98E7IBZNBATQxnA45Wej4pF
Fjxpkd05AEtHLegObtkwRmDpwmz8WiF1Q02YKozM5FR+CfctMDEudTEvERLED4XZ7OMEtTSYwE5K
CJhjjzPf1LXjIT5c/Y0GwQFHTmgf1AWFvbQrPZKWcbgSbk06+HWiPpJVWC2B1fXUS+DiEj+akleQ
6WpOv/I+xNTThd1/qi4QRGDjt4cyjH/RL5PEmUux+d/y5IJsp0dEVmFw0Ly0KT7H7n0AfL79wdhP
me5NphmELFPI+mLpm+z9pML3SMm9hkxUZEDtDMN52uDt46iwb2xPoA8sYNmURY/wHG8DgPhIBrhw
U1yMAGCEDZddW9Hau6lfl/aJkoWJliA4p3TecuHXEvu/phSS2JYkqD/1B3kPLp4L5RlTFjzDiMis
ypF7BDE6aEP+g+7+ih4l/cbylUrr2J5OyuS9quyjYWnFnyWZMfh4MbvoGbhy5y95Y0duj45rSAPa
u5aUM3RLLZn+eG96v8SBDi7Jj0ma/Q5ox/YZ+GDYLEUZKl07KLCuGyQEMwzgn+IW/glu9FB5FBEI
4OZw2ULHKp2zCcQWC8l3OUxe4OUQ8QOo8opGKwoNRZgTzv1zLfrRCZVAjrYApq5okxsPDQ+FFQlx
UcZ3k6+ZqYXar8czKup2xl/zvcFIrnzRgiLjIqSzaoAphbDDDdnV84v1iAdQvt4uWEmM8F7FbOWg
ntT4axpsxhgiVlXuGIkL+TeMThfEuvfsiVo2WghK0bs0rv1P2kzfwggQiDn88kTisLHNdZwV3OjW
qALEx6MY0yJNqBKcgZn+mhemZ6ULfA2kqaWAMIh9LBSq4Lo9jCkc3tsmMQRpifo80REWdk/ACrmH
fZN3B1Erv6F/NKoexqwMqr37yMyVzMWuFZFGA05vMRVdwAw1k5x1eCCSNqIoPsZhZqBFqfR1AE5v
aSyun6YGH1NfgY/B1qpngZ6M8ykrNnNCopvTjLT86xc/sE3xJ+yajaNWrsJFSWYtl2SQ0IOgXKtJ
irUs0egrSMhXpgPDSxJdS0tgg+1KiUVpeLxp8DN6DzUC8KDsWA9JMep0W4DkVwpnt3sUlfVeldt8
ts0y8a/NYOnt83ezQ0sPnvWRBVi3Jt0jgfSzSSWA6WpPnZhpVz+E1uJY2eQjhszBxSr9GEsfLhiz
3ocMWleVhnewxRRekZRYPjibsC3GbK1aJ4d+ixd1jVkuIRkTdgzK1HjkBK3IUkXq/TH7pBAeJ5Ri
1P4M2zXjizFrWNq+p7KRB5BrNH1EeozTpYT4YVqd6aQSmrthISdQyE265Xo8gUPBHelVZ5KIbodF
eBXK6YLyWzU18v7TTzSd4/o1G6kiGCP0w0+0/FkYRTW88aIeyfVM1E51CKayLNIc0Orzh6U8Fcfs
lLab/S4LXUEgo1JhRuG5q1IaE3xfVDqcK8+qcwcg+2211e7dZrO02zM+ET1npY3JoM4Dkes+0H88
5CniQC2OqkFcLlnW1b5UAvH6fuIBkWGHi2y14KAC2lVfd6SlhizeQF3eCECULUjgXJVylYOljlcY
xU/QoGtfpBF/vzYXGtUp+LU44jo16f2lj/nmcgBMFm1gt2N6Wuhs5epeAkLJRFQbbWFTQ1ZQUPKs
Gw/2ZT1eew1c6asBA+916S8UINl55pKq9Qxp6M1q9rUKf3/n/J6anzJs7Mo/yGPOfgtijaZDJ84h
aNvEnKc8wP+J/d/B8MKb7bbL78M9f0hhhXllD6PG2S1D0JGdxHWDZIVSpiVaBUi8PsyT+bvViUBJ
e78q9heYavEAvAJ1vqIxbmd47K/pxCjywx4xAzwADbmC697L9xy8tAEJQyweKFWto/7ilViN/wkg
UX2tw3URvA0ARn6ZZWENR5j+de39RfghQj9dSz6hfXw1JfERH8FtN/HEdT8Bj910FXxnMbooRn76
woJOMVxCJcWgTviM44Rj+Fbm4MNslYuT7KRclDbcgLPnUyk2KJPNiVPyf6A8EMy2EeHeIX9WpikK
/S/ZwANk9u5QBRnkZk0CZ/N8O2rhf/gnw3OMJezmVPqtqEw+Ogh8GxH4yb3ZtutuTsh3ASfXZY7H
yo8G22eNz8xbMDgW2wF3kYQgbVojIeQPXplQ/YRKLoc6373jT8fE2/PToieUioEDthc6jsR00zTB
+r0qNWQ2JM1h60taakNXdB1JIFA+Cve6KQMbwcaEcMjJxgluaX5ls8BCCriequmUJm4co8UlRpSL
N0aFredjxU6Jz0EgRo9IymokKg4Xhc6/JKF8KEv6JXvKJ73HyL/4JmZXrK4Haceg88mDATt76Uci
3OAWkMIVcx9BkirsNHgwkMShZ+WViZofLQ3dEbgtiA6Jybu54BGHbdrz4hzcAQ1ZSEDHzVFl5Acx
WweHyQ9J1OAn47HOPi4iDLpWPlqianTffltEIYsjUI6nDsXn1mWL2gZDffKdY75N+wj5b++4lrYC
/IwEjgyf5TDjjlzma8vbib8Tfi0Sb0AKU/AVNUL/Np61+joJEBNah/4OI9xCCVX4oiH6DUa8xty9
CDt2Qx+dF922KhSOMW1F5Y7UI+xXCuHs3+tZAfsq459U4jRSZr4E9al67DpGhn+fbqUEZA6v7aT6
hK4GgwryO3dbqBSVjZg+pK6IIjDE+QcNKlLO7J+6H3yQeSnxXcspWNmEft2cWG8FWurWLt9zrnul
lC0U3g+FoGvoxyllpGqgG5gBbE+BFg6bi6ZLzixwdt8XaQT5qX6WGb0/AXFs1WRJ71uYNgdix5VL
1ZpyxswjMoqJD3QpxpYbUqpkwo6xDWKb0eaH1sMT0fZ0MqWMTZJERKavcSoXHeEWVLQLqY2ZDDI7
5iVlDctLB8DIYCTj1XEuO3WGQEckiA1NtuowMcayC5AOR16u8jfZyeEppuFkSP9+63kDO/R5iRxg
8Uo7ryCpYPjpeAUFSaQYVY6F5x8aVk9notPQs+fBeFglkP6BmJajRYuz/weTBe+JII3sgGpK5X4Q
IrsLkQNrXtQ9DDadw/JJ8VkCgpGhabsHmql7xjRdBbiWK0Zc1+WsV9ZrqnkncWT4Z3zARq5JBRr/
qahR/d4r9wBy0NN5MX1UjPH2AGgfgP/kXjhouvcwfX7NpEv3K3VmRmEbzzpG72Bg2Ai8TOMfp/Pz
15skUEVWewKBRKevIghdUqcM9ciOjXqJfFaX53267WHTg3xD0+EgWgN5IsJ9Vm+oP+87HVHS0zAw
Q1V9VChMTtFqu5XQOYD593sYOs4merNP90QlWAKYATYDWGIS2CP51yJqH/QoC13CC1RIxCUpze0w
1D8lHGbkA3RNxwPlqZWsEHcZReBfeuFOe5XisqdIM0UpS4zbhpgxBwCKBL6qeQwLgmjlROMKriWA
RFejWWnXcROjgYuZWEaE+/EBTHeWV15RMS7m42TvZq2phpNuPISeitRJfVKNfStR5gLeDxLK3CXy
rcaYiqsKFMyCIkOQkg89KQ0LykdRPyN35PkdnpY5HwxH3JJcj5tagFqlLWcDJ12BEc4c6x/dBd0Y
gy1l3EwQNqjg8UswXkYg5E57V8RRzfqcX/y7D79LBjRfKT2pRzHqQJNBRSUnwg+nYGGe8ZH2s6bW
y6x+Uni2HqMa2J+U9u3xvSXYUQTcMw1gkuSe2rX2SqpRTB68lxS99MrlAmw5D6JOI7gvVoLQVJhi
OQ6hzIFxwp+adygvmu7Zs7Gyew/YryOXUKB5ObeRDyTMHIdQ039klI1oY9fCLTXAItFwFoSzDPNF
giow9I2oLwjHhUqrQHpyvZB9xEXph2rt6m26rTEceHnqpn/XMBaZXGjXbmSP+ECkf2QAN/C9/KVu
TBl1q1R+5CsnKCvZHRWywYa4Lngm9FTjBCUIslFXwkONMMOppNl/4DIK7s109gX1RK524bVQKL2L
GzP76jRygVz07axvslRKaiQyXqWy2S/8F8z1u4kdpnDkdZrMQVvRkq3VyoGH+rjl0HrCWs22vMP5
tmS1IBXDxu4DKza5WQxobepOu6OofM7vxMN+MQkynF+m0PoihJDVe8SxbeQJiL5Mg1schTbwoqdE
Gdr9X9gDEwa+D0ir4Tau49YP8cumNO/GTFCbL31kCZ6eRQbtHEvvh3yg3gCzvMUTV78PHHQaDjsV
j+8eGBrDsxcLscESbL09tbmkO8xz14TiUfI2mY7kzVsxZxfOQjK6Rd+iQTYODtWVqxSmx6XY+puP
KY/dujHXZJETz58rKbUf12ES351x2n/1ZmQgH5sbvHMe7xQS9mvF/I4YNyar63ewoe0c6UgSjwcS
wDU+bYDiPAYN4ygZpNm70WRL0F/NNpzqkPeZvux7t9s6D9/PxU5s0+0WKJu6bM1E9AHjVLBBEs5+
D4dd9j6iYd8bJBWbtoxkFVLZIsxfvIcZAkN+wupqbqCP/BLCQD0wc5GJibTvKnyvqwfKF3h4fVA8
q1VFPs8Kz1tZQOARK20RIZLa15aT20LHJ8Jr14ZSRXh2PvsB3SwxrfyylS3wHjGC/fFT9k/WyLNQ
7PMMGQaN7wiE7OGeJLTvlvqtikG7niMxHfLJsOHoZJYBp8SIz2PVHokqp+p21ZCz0pZM0GKNJ9Bo
0nBjS6Cgky3La7h5onQjfH8xELreixaBT6oeLQPhYgmWImDjf+7JCOijonmP6UJYUsBHd7ptj7lT
Wwhc5ykQRIPQUPTuoDGw4L02w8yyR+Qj9OSyr8vN0IEaFu0wWTdIgLY3998GSj4urrR+lfPCbazL
Uf59/i5VWqZVqYgWFb/UlASmnLfVwRBuIEgFyeWYw2IIDLF4KkaaDGX/HS6HggqTTKVrko/bAa6H
AkT+Kh7jiBIoYrlf7GT53aVTgWrZxXAO/8pY9rvNneHQqzckqF0a4/KSqZFBy26P2FyRw9LJ0RC8
kE0+ify2TLEInQ6aNxcsO0Gwjaz1okOlw6XZUm/65KYwYGMXhJ6VFDbpdzTmXcAwarr4pUHc2vz4
SMrZys8OZxYjSceOtdg0/BH56qz1cFi5RI03hm45K3K7h/DD40FknweFw1ge6BQZaKkF3zHmHXqj
bNvTpPnXgx2WOpxCeKBObDFCQ9e4Us+knzFIb+Mko6myS+dJtsE0XeUSYCa0Hy3ZBt6uWumyGDpo
i3bLMd8RJeFIHSld0tPXnYV4R6IzaNyRAOkrLjiAL7nznqh8p5PL7UEUagtZO3GydWZuroRUZYN0
Pf3ur1BQHZrN/yxW+veWvc6yfYKsUn82R7MGqCneQpXqKGFenewadWTrMw/KigVF472V+llL4SmY
ByJDKT42wYcp0GvfPKxD4ikgNFcO/1Zggy+JC3j0NvKwkJcZ/5GbGhSv5nFTg1IYzyh4Xsa3qRLq
uyK30JpkIOktahFv0WQ0LswQd2yYsceRVXkeDX1r9uMj954kdFY6EV92Zt98y+8Guj2AwJfdeWtQ
zOtSrBGdUbDAMcOe64xkJMKEywNg6Wja8Bg+IuSGcWMOhr8qH25eFHuxmgRj3gTmbMB5uG4NffGY
d6yFoQ7B1+kUo6MwOTNbvQveL6V/YJe7hNyXg2oBcLj3f5SolA0vJZHeRBZvkOFmiCDAGMFqzzPn
ptcQGAQmp5c078wL0BMiNALdgTY8xEQ5cODj2E9l/dj7Vt8iW/dUBHz0RQjXlHTL0SxhGNDWg61C
vXA6yhT1m/HGzeg0SKugYOg4UwOTpC+9UkTh5ka6sNO0YP5/W4iRKQCnScfF/mzYLxFDm52FqsLm
GS1Qcw8jEZbjnuUineHzmFmqldE7ty9ZLpbJsCt91b9mBWNh4R9qjhCeCTozCPUF5dWmuhuwE0Oh
dYg8gjDxLVaqNt49W6B3efw8sVtpdNOEppvNqHayu6+ZXuWlruxMdfjA6PoEzGpJGxVQdFNdfAwY
kFmjCobPNuyIjIAb9N1gTu2xbFFJ/G3GYwBagdjvt99iQsKBlDscRn5IMlp5cuJkbBrOUJF11WvR
aMk5n8h03Ubjgv5GJTx10D0aNGmwDkwJ+a0Ht/wp9KGip2zH3tRJVxiEInuh5e7JlPpD+urV64HM
XVqTxk/Bx99WtjkPlVJvq5/dE0GPnDX4hMgBMlOU7fr5+mcny6s69CXcaub4U0gw2MNyuAxWUhIZ
YrQU0pVSVswTpP2+0f4rQVoESN+obOyZfXinoBUar1UEIiHOhVI1pvwNrqAPLEHwzprPHJqz/z2B
hjzUY6TKSu8uDwT9TSj3Q5L2o8uG+UzeVtpTZLaVyrAcl4L7SI28sT+fq8syeeHLWwHN5cKGH5OO
GzhAIC7QpdksCeUH5A4+qQIHiVMb1QqZXbJNIKT74rjJsE3ym7WcS2ySt67YilaxXAIxm56uP1X1
NITYLqkgn2cpKi5I0+M3qWo0MUbllRktShlAz7oVE1hFTAp8Z759hAmScXtfWOjF7L5DB6dQDCeB
sPdcze8gdU6zySqHMeMbf/fkciqg87JdIFE+67EhLvjBUmsudubGZV+A/QuBH6G3qltZZ3tz16Aw
6IUvUu4XrSB8YYYDIdutPhkJGzvUU4A/sUx1FzPa0vuEV83YscbE4VJdEjbq62OUv48HNdH0p+Mz
zAbsrhruugpWWW8YQHZ/IgytsyJl42IRaEz95hRzMpWxhM7jeb/gBDZvgUZMxFDa6gbybk55VSne
Beq/OjLchMzZRDKtrIz8KDF3556/JOp035q3TuX7ioL3/QIY5ZyqOjIWzq2ZTBGJjQKxyrb+UQXf
HiScFu+Kk7NxtOoAkL/ld2bLCSL4ISw81DbVPNgDwUNNjOrSo+ELVphN/xFj72I3SH9CQp+MVQ0I
ELVFJaHbGigf3E+Lf/mBTt8xk+VdQy3R8EhHNrr2vl8dtMMPftXng0xk9EzqxtQQ4b5PA1/UBr0q
ovPr1CS2/gJu66lqXi2lu3wIB5af6lJceOnA3UyCCQ0boxHOCOzeAFNJw2Ian/7SxOoND/6+Fyzj
uo3VI59PTtHnn2WtbwuQvmsgAeEbalJzQKRsExhJZAlGWqsCLJgiHAhH+ERQR3oKJFfKqvHHm1RG
sEN1Tbi3nxApJ0WY7JDQeNbla1lY8bg/DbxTWLN4zjaKdyEzw+gORDAEGKoX2NC4Vvt4ILVpatyd
PDoBQaXn077MrIbKWgR8B1ejNHewVTuvK1uGZ8/qZj1YBG7oXWcfuEQHo7kOV0fI74TPFcbiDBMv
27E7KOS74yo9vcW+SDOPZq96eKlwPExdndTSjmRrRQwlo3mq7ief13VX5tZC7MTl5CVcLDoNOw8s
BRi3sIK3FMTFpWUEDo8rSYa2uHZnIZqisk4p5ioIx/V5a641UQ2okzXilv0SG1CPAI2HqnUoIzxg
Pac7RENnXCnEhXw+Ny9aG48Q8+nbrZT+Aj+JgCYtgUvlm2MEWqjk9PsGBl/+/s5zlV7JeDxcBgQ3
QxJu6Cq5AgIZ3KZJWmaQiSVtjpwkmyoCflXf2I14oVzmczjlAa/41wzZkRVdRvjGX/z2tojE/MzK
L+R8R4uMLODs2rnXX7QdX80svJ7vm4kUO0TDH1TuQwNBp93nDdHe07vsiTmtVRSp95FTGwccS6fY
A14R/2DmuIL7Us7jU/s9NKQeOghMy/f/4qbaXlzNYNkLeeLEs6gIRbykJbhXKEq0tznok5Eaa+UK
a1MTKnusJN0DL20EWV/oEyvRirzyxOUIFNtfyhU02UIjplAzsWiZ12HZeL5MFZ9XZtB6w1Du39it
/57ZtP001Q9g0JauT0odHU4Iq20bm1jGPqp6JEvq1UhA7RF0mVSV02RZ7cABW9dK7l7MqoKrOKCH
XBCBZdKWBsc7Q+V/aE9zFBgE7/XHrKNkEphQ5zcwKHM8PN7Ci2geR0c/Ysfhe9DRVn2KN3uSjqTR
Mf4rvDSo8oAR1dUFUWvo/I+gfhyMRuKCCYHxY7+9uRYA5uOkxSqmkwyKP38xLCMu73z7PanVSg4J
0tCPDX8rGkoZP1Zczm/Ooz6enlnU5pjJX2HJs6jCSugeaZJhUReop842j7EAm9i3vh+bim2AWu8C
k2oYEheN/H0loG1RK0vWjy8hkhMoY3L2EF61phfwP9N+m71/Yv2y52CLhUAQXWE2ga0OQCVbw/Kd
2t2jZfBNF3eCGMHs6FvDIyFHtxbs/bDP7JYECgDtLhGKodn18Nlfoiv4MeC5dibeNXigk5HTFYnx
H7TvU8PBX1wTgdKslx4m7dX/v2UBCCtpqb0IbLkDjZMwmivGFSvCs8vPqwfo6eTo3CPuDMwiWvf7
2n0fJIRoX7bYQRHmMawNjQ+xlH/sPYwvZcY4kpuZ+XP4ijlvGnQTsF/ivx5+sD4xLNTnaUxHAi6/
p8yCsJOY1nJRWwoWMW5WDrTMnmjf+jhRXmcAYIiRlG08oGGbupFTqFj/4BYmDYBzIwGgtoHbXiS7
yWPfJsCXqhCebolVqpScN+0vorU0MQ6D/VI/ouAPuRPFNEsq85X/5m2vSM/9+dv7a42WhRTwchAx
fd/x+tjDGoHQR7825/iqfpIhW9OgKjhcUt3jO5ZlKgQmTMOoFkpsLViteZnPCL16veKUr3ZGL4mU
tCLjNhPooJhpdrqid6y3Fo0b8774sZzWKLlRFJ34XFJeUeq8aWd5YSA8cJQvg5RwN8oMrWWc4ITL
kurxtizqzc0/saPpxogPYqNBx7VfWwuOVu0x0FRk2rn8LnSMjFFvlsNtP+1CqYV41iiF0SnsiBuw
5eKrbthVVqCNxFaxcG7iPALiuCbntt/g6vbnXjtp6J0hkBg5dD1edGfeWu5iKjmo5aKSb6sNvCkj
Feq/KbiD08oPTSy7uR7vuXagGjINkg6GrmmSptf+k0owqvUV5zkBk3fa1SM6HFVr+IsDvUkAx1Y3
zSrRaQmtLBi1NQar912HC7NBnveyi99E53CydTuW3J2lNy3N2yMBs4634JrOjtNzdUyBmUFSZr3u
52pq3zx7Mkg25VRorD0w/AEaJJ20WKxdxX8vBH8taSUiQgiV+vuZ8p0EQvNVbpfBxeeWnAWIBv8b
lMto9ZW+tU8jr8gCWjL6ybiYC32fYmLlYiILuBN+LNXrpupjh8b4Q1vyVZDG1jSQbT2dHPrUGwxS
osoWx3/4WCSNQzJReINX6fp/GizN0VTb3u17nXKmujYmSsfI4RaYk6N4k/XomSk94+My0reiYvPX
xerE4qwmEdvfmbncFH+tRyQHG+B5/Aby5fjv+NpuPf7El3Kt3gjV6L4vywKB0gILOw/s2Zxjorbd
7+QtojX4yvqeQjl52zp8njkZ91HgzLRy/cZYMaB1IH83qyruCrpPUaw+GDajWNSOcNHIFxwd5FQx
h0tgK8pvBNfesU1Clt6XcOXl2bgAsOJDA2Dlp6AAFs6XXP9zMF4cqzCIju5HBJdtikEHKKaStBuK
+0TIFMca6d6oXURTqwV++cLUUOGg8Bo8aJorHPGHO98h8a3Do6nX3G/fxebxIxuwdzNfv6SQHwZo
iuWVEfw8A+9G06PhNOl90QOp7CIR6jMd681PsSRJnsdIjlO7NYht/n6AZsFkKcsawYgP2WXwNkaU
goU8fQMOc5DopZyJw6RD6Rlz+gzDIjg6vL6NU87WmvYOVfYwHW1mQIXnYNwRr5tUvL14qx4zpCP1
2dDYBf0MVLT2thsW7h28BoJxvBNex6jTN7N4Hos78njqhSe95drWJ98B2ZvVYwJXf2SRJWyNlMII
fhOxK2R7B02W4udf1Bt7FcP6N0CXS3iotqigry9rlY4Hzdga4PzrZS08PNX5XgUwmDJTlFgHP+Bl
xq2Reiky4/jhFEJDULDx3TfPn7nA/pEwaYxft2FBsXgLv59eKfRBP3Ua7bKlv+hGliuYr1tWUfI+
SlTj0li856JJQva7cJomRI3UcvnVZpXbxeFWJikG2g6Lke1RZFWSGJBHfZLJk6i+uO8V2gTKNNs6
0VjR+OgEAzk4NBHkRiNpdDZEMLCBYfLCYnwp5Viky20Xs+xAUoLmfynIx7vAw6UjeeFQG9H9lOSV
hDOfRej8BKUyJVeVek8PxNHm9MaFfAtfzX9es/A4QZ0IqFRLIZE5fz5aN+sjFFST+QR8MCudc7Ia
+4+HOkOhMnBMYBhQy/9y8z+FrMoYmo3kAv3WwYYNtIt+M1jI0R7JPUkFefM8wEu5dpsTQ6j9nIUo
9umTFVROXwCATEtbAl5nZ1zh2Qb23KwHGh7oT6P/heR4poUW9ClA459kHi0V81333kRLi98xg6uZ
wkmCulDfH1dF50s2oV85IicuCZ4s/QyZBLj0c/2x5JO4sYuJH7PhSIzezZo43A6oF0AzNzBvKAHu
8IS+iqRpBPOA7Vjdxnr7HaJGaKEpcWxMx68oT0Tvwv7ImVpFU8pPrIfTcHz2dzvhhyZqZL7Q1LjV
kFOzevBKZsk2FskYBRnllVJteRATdDnYTQdT/ise62/tR83hFW+m5iC0CIzfcHwv/GG0OblSdH5R
PV1O1Vx+JdUr32UPaWrYQwIP0EfPWXe6DYsFIdtRtVld0n65ROp4Eqb38Z5jKFHFEQv0IgZ4DuZp
RnxKNGEsWcOHPgSouNBsxMln+xTqrEJbtcGLipIviYVqXce7fRUdUCEgmhD4Fv2QgpskFPG65j2A
J2ZJQL3vg19RZlTiFaWbeKTi3wUj/pn3dOX6O68p16q/uhnkxstomfp87jqw5sFK/RkJFXnIXwHd
ZrH3Np7QbBCeiW+OgOQcO0gecMJDLQjHwX/yxrx5LTCoeVik0fkXjccQp7hebdSDSr9xhbTwQt8l
8Yysr/A8pQYjF1ag+lKbk+J/+8oFTzap6k9LkkpKGURQmLeMZU8m8gJaE65qJvBWqvXc1uuT1Md5
qbtVlyGNIzAtq3rFd6J7GuY9xiAUuA+/5v01GxywwD6NidOVbFT64xViuG7Iv/c+cdKAXb7sFYEH
hDGVnz9PrDS8nKClnaaS6Pm3KYvfmUpN0TDL35KquOahHhlzRAOeqrm4FC7fxtwvAFDzzNGkqr1m
0StFLbxSkz6CJKnBQQBPTkEbwuYFdxxlLvv3O2kfnAMR/SiXXqLRm1NAYIzhbQQ/nfbWEBDxF0TA
jYiQEBXLF/rs1BhIwON0drzHXEXhmjaltSFEmolwBgEseq10FIi2ysVMtaf2idJyApg6X+OPpoKr
WV6cRZg/RMPqj6Nzj+SCOUY0Fts0unBEh86TEvrNj39M/N7jD5d8uXeP/QwtWiKmbzKKxeWuPWfa
0UQmTTARtmWqWajQ4EKQfQvL0IfjsNdwLTrBSxaMuDbno8kZZshEth1fS4MwVOB0YcPbA2UXl4p0
lfy+4UjsG6OqXRBChi++i9T2Pw==
`protect end_protected
