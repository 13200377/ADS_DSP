-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
mraLKAWKGzO/3F6RLPvvsHG/C8TrbkjsoidUQuu1ef598JoW96TgVTOYJ5axvO7GvMTLwZnzfD41
PwjCdbAfM/jCBT6RA3GJ1p7sUn1S7rOXgmlhIim0LErR8QwI9xn6rw/Cu4Am7wSRNY5bO00jFMp8
kCOLJeaOGadY5FKb7xusXdVjD02iafxibCOSKVtMiX7L1zlf33uDu8+KwbCpNoKzxGCJiT3gX0jL
beVoJlz1w6DYZDZXluXTZiNiTeCMXo1DxIXglyMHQTeaO4MmM/+OKYpro6zs6PjxOImk1qrgoyVf
NlYXcE/zHcFg8bdk8JPBo/PFQBns+g58Z4CCYw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35616)
`protect data_block
P7C84Kcc3akbC45Va8QOmfqRFbx9wrdtlMzYOn4l7YGC/Z7f4ZAGd9hLjCidc14mxKnNIfLiAVNM
VeyVYHQmjcEVzIAuZE2a8yTeIU9ZMSnp2W/nuh6jsu8tT9nLjbtCXC9C0a4/jMxeuULIoeekEWBl
0mL+XdRpIWA7/shBrdSNTuJrO8cB3N8R0ikXh6RNXESZz6zARMRj+J7Ez/2l46dHRyw9lxqgfwgj
Pdgj4rLUlGohr48/6ZbnENUuygN8MRtxW5AeorwAEfmLSMyHl0ZWH4nLAVrU0bvl/1Z48Tv7vMiz
tuexIBLjIxSxLRWjzEt26c23K9ojrK5j4o/repQa9K0g79r8JEhi/Z7UldaRgjhbJcm+NxjWCBQp
MLBXfXiefWlpdc1SYZwfV5H3ppfVpDD+9sBpGplat5Kf9h2kV4Cy1/Mz883EKGwINjyc5ymtL/OK
UKrExa7uCAKDb0BdmwpUadpMzV8w9VSiK9d2grY1bDrlFaiRNzK5GsHR+DPDwZRZuxqgM38KV4sU
ZI/0CVhlkO6aAm4/KRbCqPkpDjNDn6ggQ7Nm6z/AA3W+BxEogxrsIkp+gWdW3ev7F1Cx38VYlKFa
I99pqMuDcwH0F+OsVjaZUvhgPhizKXoMBWS6vjtDVc2sUCRdWNoABPHTRRSUSA7ayCgkHvRnFwwa
araeK6G9XTgmuJ0TO+LFNG8P2DHRe6YSQN49/q9mV0MXSVgn/5vxskjQfP94P8PvtArE4Y7I66yU
dnbkSL1cPLQNMR4iHDMh0c0adSODfmKs4ZlUI0VB84NT5Shk5Nl8MTusCJu/SccE/DzhQ3P0lkU/
FGuTcrhtYZ/KM3VS8SgeiIqwSPpc6LdPhMiXkRs3Gx/mMCg71IUW+EsvaFcG74Li0MFdU1/yZTmU
Hms17TaSAdZc2e+07fNM6K5u/s3TzgYs4/H1s84ybeW0bFOa/AB+ItDqY32yd4DVJNXcB4ZG9bub
MMxyOABk3jdyILvA9q25zL0lfdyMWkhC/1YZVNf6uEXRUvLRdZAbxOZjTBo6XBWmQlYvN7s6zZm4
/B9HWaFbPXvbXI7XpIdLRIRK7jesLRP7GVApheV/xe3bFU+QwIZXEQpp2v7Lj8Y1gGRtGijueTV4
9bbQkQRhAhCg9qnILtcOtCLq+JSq92RcVTfiKhvKwY2OQuecoIcAu7MtVlxXMnBDyPvoXb9CT8lz
iJegJhminqcZGvvBzB3PcOMVwZfttMIrGJlCqjMs8TLG5o7dK29njaEvNr4GK1x9fK4GXgTnov9p
i6VCRXIZ9ZxUA+eYL3/VegMVgmTYwdjMcEa//NCSouslZAJd/qSsI5/3vMQZTHGSQK9QGq+VsIRf
+IezxulRVFbBx8CvhL+Z5mb7TF324woso7Uwi4aQqMNQXEMEeB0iKaweFOqx4b9m9mR3SDjb6J9P
d056Z3f8e9+UYe/pekySr+8sDgWxmrNeIIjxDvVIwCIPrn4WiNAAsx5UaLPv7U/mYAzJMrvUp4Nf
fZawtO0BdERDGGud/epyDP34p/JEeG3JDRjhrD4Aggcn6olvlju3wIa/Wsy8J9RuIV7/FH02dlfC
G1YONQOeAd+kHp2UGTG9gnxx2Yx+MwWzD/dKwi7Mu/QsC1H3cBuzbvTh5TpFq4gnTz0meT3GIL0u
wmbthDfQWfREtHxmFCWDtBBdsJvn91yXl0XKdRd2pKJ9d8hM4cl2AMK9NHHpxb52VAk4ZC3NoVJ2
P8h26qCJG+JocNd5A3WulsQ3Lh6Y4MbYANLw1srHvQpleC7ArpNsAr2gSZ9FZkSB78r/pszc3i0K
Yot8XD8k7pzrCKmO8Av6f+vFPWe8t97N/pHfNgOn1/BJqbH40ydkHoUNmMwJ+bibjSGsdfBZV7X7
3vNicfyS5AlzEp0jMx0YAaWyEp/ryk+yH3K0zzuOp52v15iXBUGUXMsnndQ69WsCwfoBG+F1gr/Q
OstpnkStTimwI0pbtsFkCRsXJ5Q0SFsrTA8IJPxNXvH4T4LWT3SNSt70IIRWiP4U2dFWSWm0yNyl
NTTE2FQSEDFQf3FicbDSMIQVC1eg/DBeqAAujXPtL7BA13nZ64kzfHeIsUtmQg8BMhqHsTEHpU+B
gK+x8LaITutAMtwk9vGjcsKadLrRYZvxY2qCm4tBVdn1WsU9oMtJHMDC2oQC5HdNdNf+2jtN9Nyn
2Jm7cyq7ldLw1HA9rvWJK00P72vpf9SrsxOMn0zOM15vs79+Q48g5Ity9j27OyxsW8oTcNjW12BC
R9iElNPPJBqWrETqUQEuY5sqlUdfdOh5E6qLriNGxiOVFzh75Q2ubee+p0j1qhEjBUuW+YmiwPXT
g0qIp6T3MjpNiTb120Nm+Ui3v8Ioh5Ca/bqX8IH5WM6cpIahd4WL/3+kWRrd1r4FA8PQqVyajk0t
w8uHfBri8Xd0e2XUTRVlyWhvyilxYrFWA2WuaIrGHZ3pPlVLmvaSfRmmiK3R63NU7A/MJCHeoUeI
WmbVOoCExcfMgtv/e87WPx1IyHOUnYBEVLYluMRZmECI49iK4UXFEGvoSJ3WZrZi+ZWaNhFAV/rS
6Jus62d8sRs4NqTCk0jpyse5znz7QcpgxRkJIMDnPJaNZFGlZgB41l+KmE4fV7ZzcWdNwmMNcDDH
dxg+wBEYyIIgXl5ldwLb7nWLER0BZAeyoiN+w/rmVpoq143uiD2l0wEPDjnHo7DNGrZUjjmEeVHh
kDoPnsb/kRfB/o3tQrEJeyUWOqmBMB3FUhQubmRq8pNu2ucAthdcCKHowC2emCSOTE/HIas8D+/R
/mYhV9pmcvEyFYH2luuprmOeMGrBhggXMC6PiD1A1oZTZoVSCtw2a049GS/LOWZeDAzQdq5e/tR9
kd6sZ5MWWVGzcz4AbjjulJNEHiYxYjsvir2um2OoBpLepU61L1izXNu1rgBs+P8o34G0CUPdjAe0
VgopK5nDIFCNeMhAHcV7snKegAKWgyOBvW8EvRxDrBMPMyhWQVmJZCRXNnQGsKlBp4OcNeS316Cd
mYzqW+VxWsNAjMyIWPzY8UWYxk+TN8PWNPPqC6N3fYfc9r/6TWDn7jDE0ybFp6HEKFTg7Tm0X198
CvHLc9WLGy4jJmlbcyqeKJzLRBgXG6vKhfeFGHXZNP+sjh5twl+bBR6W1TnbzvVoKqQK6Zcg8RWF
WHyKGnti/+Ue/mMpe4fitjJsiWll2RTcYaHQvcCnsK3sj7+K22b/ImPB/aiHPQKswDezyDdLMbGr
C7pvNzZqF3Ya7y6bDRtoaJcQiSOoPwEEtk0+IT1fxXrnEks7/IBeymERfS0qBU4gNyMiJel9QWzU
LU+mPD/nkFWSR4MoB1gRzHVgUSNYbjLeqKhaQsNh2kLOwjU3aEAfDEDknIYyJab2p8D1z0Pljg+o
C7nMoaKIqA4/qbM6qzRF6TgWFe3jGuDyU5ciMAX9Ck9TdYOS4eagy1YDc6AYRjsWrcz5Yr/ch/d6
B/TVndUhHNK46GlhVG+nq6HB0k2gMD2XG36DjgxRtsdGJicgYFpx0Oed5vAZRI15Ttu2uryK4r9m
imT4kmi3y7tBa7AVjOypSg/uWAB4mMEefX3F5lKG1ZDHEtx0G9FWTq+hrSQZcQlsjy7qVhSQYgqw
ZqJ8eVh5DIeB8gvlYBEyfnJiijkdJRasB7i4YQtX9/sQkJufo7ZQlVvmkuzcvLOKKBqSgvOJu09B
sWVqGJCK3TFy+716sY1v+nS/e0Lxvs3OeocOI1gxEpsgual8wIoYMdVyOZJMMMMxuWnk36RQoy8U
cxMMqAuKbUdDJv3G/OtEK8r5HdrET/FLirxkyqdPHdEThXKiSWEGLt+L1XNFQyq8rrbtAYu1rU2s
5Y74fGQt19Zj3FJe7k2nOZrtvU6srSnMLygm40iCPLvTDHggEqByTGoBodMDsEDcSZjB0818t+SI
13Da0q64W2hA9KfQxTYytFkfIlLo0pMGOwkBi6wa9WqIDiza6ZWEQPw8LmS1lzQzfhvKXMFOo1xw
IHxqM6+2F/NsBmD8PAPiORnZ3DK8HPWlR4KvyVOg+J6uc7QrNdH6mB+WHuFiJQmzB+fSOORqiS6p
Id2MGFdWyGt4i47lIVVm3WMmVovUwxCm3uJQV3C3xVIhyJcx2vd5kgr9ZGqy499hrh89XiVgOjiM
egAxJkqQzvast6flfY+DtYHRrgIzC0rI48LB51pnjtlPOylJ5Jdbe+0oAsEVAUNi3g6KHL0duc0b
U61R7L7PJ7Qfezt72416d+K7tWaVcV7n7hyLP2n/ghvRImdDAbkUPWncCGL/jusKTDrwmMwI0s3h
d/wle9wn36oBfi63U4tvaPaNRewQbK1/KG+KmJ+f8cZK8iS8MLQFQNHynlFfa+rymnUsVZmveHmk
I7oP6Ycreu5i9fJRSgxTWlbfgZZmBKmOEhf1gKpFiNyZfa1tya9gLk+MGUIno7vZGqijNsBaJJn8
K+jcjGXHUjvEk0Wq0EctvcrxGmBNSGQ8ngwhi1kRcAj2bbNDtLjPq6OlfMWBGgMvXWxudw9J2HXp
2bd6q/+BUTF6BnrsKzIC/MPp8os34CaGyjQkjX+mM+0d5X3nqzoDL91+UAJmLqv9OVjnI2dvVWCt
K+4pJEeOCdX9NwaQEYpCbxHol8j11hFIaDxAuVwfrWLqgPl1kWbLPgWknV0ZR6QtG2/HYrwmr225
PYyNqECtfKf/wOSCisUfPBKA6c77d2Gm6L5uvoXKWfNAj1y6axim1xSNLtO5MtMS7B61ouIRm6Gn
FZkm3vw81JFNuhAnaWW2j8/vd3PGE/VYf91ia0KNfBOobpF7WgPMZTzaB9vW9qxVwGeGGF6MqGzt
n5x7TCCgLb1L8p7RaQe8qRwYaghbG9kK9fcPwyPlrLfkeZvN+mU1MOqVXov+liGmGljDXA4vv1yb
9aWbNeaRZYPFqud+37W/e9LQKQwyLFSpa3sL8qx7ixtYTqvbu5MTwKd9oz7cUslwrETZazVL+ZP0
dG+8muWYGPombiKhjaxsVNEY1/cBWVWm97dVh08mYc2e+uIqbSt+iplHHkcIHf8u/rzGUNZqFt0f
5Y3dVn7srRzegA/U5bDlRPHLCwuUIZa1LWrhVUZAT0y7rx5QJBLS5CHi17ma0/GQT82jFBah/btt
6MbHKqGkclludQPv1m93sSAf9vm4ToqC59J4UdOlA5k3j+/rMsfew8USM92aVqZBzk+qN8bdGmbQ
PR54JjJ8aSiw79IVTVr9ouywp+LI2rizXmNktqv8UfzSoIAValYHEvR9Hw8JQmbJ5QeSief/+g3k
8Lb9TmJkkRFWjE0G7UrYwhtKT9jSCToo2N3Rlm0j9HZw0vRWsnS0EXMFOcPwY4zBB7k+HLGbimXq
Vp2gdg6uXx6gbEO9qWywvhJjUn+PK4pxHlTRwgOCFyIMVj+s1crnQzcpuDxWpM8tZmLfgZS38iqJ
1GE0hmItHWuuudm9A+Jv3Fof9WQLpIWNCubdLVs3icU8IM+fX28p9qxJtWLScJPZs4wBk5d0Gt/2
R0nJolNVRGNuiJI84qDUYIHSP0FawVfYq5YmLaBJ98gKr2N6Z24+0kjQ5O24KocSIRY9Grxuze1i
H6DDf/7MnCnV5oJGMGDzH5o/fdrhqnkrU0iw3ORFApfP6Ydz8tZSOF3LvlKZIDgj+aQrioZv2s+n
hCN2pDGZ7qlS/ZL1wcQjq8tPr4sVv5T5yW/G4QZjILwDFft6fr/KINYvQ5Vp4vf7hFmh5HpqrogN
Lv07FON+K+ztxadzYp2Mvz8/tgcpgptBe5c+4G88lMAf68wbocC00oB+rlK7DltkW08JNTpH5bPm
JD+jFeLbhZKrDSDqP8+iDxPsN9q32sLvSNojJaBcLG4ezdcQ0hYobKRU9nPox1y8vwscN1qPl6XJ
AKT4RZptSnMhmBDvWuSDGRYNpsEqlz8Uu3YauqYs1by+/KPGWPgi0uJWFKSsjaNzzYOlX+kLo3ag
Xnt+lMDNfr0k+ssY5dWksMk3xSQslDaG+2UB9VAJa3ffktdxjoHDp7XYHD+jw5UEBFj/3YvjwaKF
VxtotBb41NcrLe5OY717AxrbLhg2GDEA/HkXV3MLugn/kvvB15y/weKp3ewYIfmZrG602sJudEam
QlQzUTJ/gPDsum+DvEL6VWVPAd4DC3ZoeoTUhjzTsvhCaIskYbZFyBbOGxvKw1cycbOnvL/VUWVA
jXvzCKJn9l/lJRBuapizIAeJVI0vQfdxYIFcPBwYeSc+1h0PoKYSVrK8ZSJ53hJqxf6r2WWfNGMf
Q61JUubmx0p71oi8ldBTw4UsIX/v11w6MwH/u2rq9j9mEj8c+V24yLFAZEvULMv/f8fpSjLOo5UG
Dt/HtszVfmM8H1t6yf9jNBvZx8JnRHh3dosg0d1kvFCKoUlms+7F52YP0CIiFoNEivH+EC8EevJf
8WiknEE7yarJaq7HbbvdFKM0eoA8Cfig6fUOAA/PA3w9OT6p7XlmOspRA+KyOdtdQNyrMEDyoSqb
IM617wKX/JYgLgFEUQU9dOZkc2NwpCwgqkVD8velBCb88rxZlSEWosdxP1w9GV+wHqmH3J6Gu+7G
/01ZstY+2aRrLV68baXt0bGSEpEdqutAjbN1bIQiOD2BcT+GYDiWfSG4kjB3ZXzYXd/HkLmNlYDc
Hrz5hS3GsbPNBk70OuvxNKdnDRfczna7TJtKVh587cHmSnf4TxLliVhoyInQoHO13toITRvvDW3K
u4PQUsoo1tBJ8NLqANrMlQ6faMnre/BjtzGfFPdAUIT2kO4owsHqGVE/9QF7SEOtN/WzylzOvt5b
yGds/G9VADNep/SmuQniDV1zxMUc8FCfRg7BIv48DyBmV9SyveF7T9nsWQgm6oJbWMGnTCtOfDOu
mpY684DZ5Lsk16Do3TbZzclbnuRb0WTkE318eZ7nGlMEBXKqSpsOnLhMGItT/7JRHZHGYHTDwv76
+okkxW3UHdNGQUlXKHLxf0fvzqQBBH9/w86oDvKuJ9iOuz/MXdjsUigQHMEVj8XZN/2oC9eDPGpU
WjL1jVjB6RclsN5KE79PCQErwAhVftACwswdj/XgrzifVoVkkaBcDNvyhAy/aH8NBT+KcS9RV3Ms
jE2xRbN1xBqFuXasKD3mqD9kxfUHrc58Rn8Map8lmabeylVrDvjSNovLQ6Vw2Sr0gOWaznNSyNEJ
OXtmxLL6cs43aBwPc7GwvG1l6NV+dfWyn49mGz6m7VDke7JMsnFRCU11lBOtVPCtUorRG/5h55q3
msWAPqcCCngg7oawAgiG2Sa25BxFuBljqVun6+A7hf178jmTsqQbaOjCkGLWE6Q6A2W6P6FcItyB
cH0gf5b602Z6ir84FMiH8Lhps7W+R64Hd7MSPDk0IDAGV9Ld1WZPo4MhFWarwp+i79ivqZ2hckga
OrrzTG8nTXR7/o9aLeFIXEoswf+dL7TxVATYlQ2XpQKP4DI+OPx1xf7W8q0JIh1ihBuVGOCEjO6f
8zpgovE7+lBfGRDqY1OWctLW8nOMF+5b3palIoj45G8wFW9k96KLaf33M/gHuI+bQ2HglSmSlg0I
U0idMae9Mwjr2xlQ+1xioocN1G4z5FXkXElT39XdoDU462/7JFRDgekvFJERG3/7g3Tll4KuRB+Z
Qo8W3k2einD0lKmrhSEtCtAmMOs3SIVq1XUjGVaiN6+11lrzBy3hb54QClNZxQM/jsGg4pc+Izxa
ceJBlBVixCBjztROWgIxduwRUFLEZds26Iq+S91GU9slzs3lWg9PMEe4r+tC2vQeRHnC28sMB7xB
JUihxWaTwkJ8PTrQZ2HwYU7MJG5a3QdeQ+i+4qnCyk794UXCqZsiYhkiQC2EoFkktawLTyNM9Wzz
PEVFnxx/EMWpQf77lYnICdsLkXHzPdnzuMOZKjq2vQuOe5cVFQ0reB6vb4/SQy2DV9YSBWdrm9Kg
Or8bhLac8mnj37L7GDQTW6YykQ7SWXPsMDOIJNAfFcRV78sVaR3R1PnydFaqQndUWgHYhFmbsZNe
02BwIG63eAlFuYrS/bAUCzOg0e6wAfNbrNQia/95HMrDTWcdb9YisSbCTGBulIiI6LDC6Qo6GYoT
Z8i7YLsf7dgEAPQsLtUnoM5VWzKSHN73EuUmIRZFvkEHVnp6+F/gDCsxumhQ6o+657bYPJfH+U+D
JZXXsafPK71uB/g0AlNm17XeRIMwyZfEus/7xKDrrEP+ms4ZzRUclMwrQ0BkL+eohCWEU7lEwOjl
VzY3uoQJe0/5TtNVIDAFCLykzTcJtjWsAdTduqCSSKVBDVQOYTq1uwhM9MTqZbFIUAjDqFY+gRJR
uvMJaqPf/zV5TDrRJKHprrEZGkIJ64jy6e+FqUTIu5SHOnQD8K5JjKKsX86XfHNOmJcyJmyC3w8+
LEoQkG976sIbg3Fx2nhUItLtTbYRL2CM/L/Vc5pZNs4z8m0UPwZpu7QoZv8iTe489kg6inXgvafQ
2ZWq1+Ayn3uYJMSGrMeM/8B5ivvHwnXmZWrMQTECsDsfKCjJPOzB6SwGv3soIfeFXydw1NLqY6jX
LIGeNjfhrc3M+zf8hGX7MamYls143NsFsaKv5paed8l4BncUYd7wD9b3/qCtINA6UCRoo7xXBkcu
y7GRA2vJmbGU+iCJu3KjNFzgWCtBW3iomQ88+mmBZmEv+AtWSIt9BsMJzsp7QvWxunmBVD1ZzrK6
D3r+ruq5Kb5pyzDVbdO38yH6XdjOHAs4TlUqrPcXidynyLoFW1NGVgRJ9rtDWsTUEtxfqL99oH/4
r1uKqiXev5WDs/IbXS5MSdEOyJxBXzOWdqfNHxhprKuo3kLtDsjnH81eAy/1Jyry12frX4D4vNQv
N/mz4Ku1WQKriZ4ZWuAVXWGVYf9LWMf3dT3TLhCU0xxZBaLcZ022lIM0vBHfADyFequUuD6JWbk0
+d7zr13nW9Z5O5geXBgTrRXvqlOPndPBGCM7fqXzM5LMmq+SoFtkfuN1C7f7p/0fN7xdaC4m3TS+
jdIglBoxZGh36inlzDGIBCcqTrAo3Kkg4c413sP43iKiBy/0O+qDdVri5ZOdEhzCKbzuaTGl6MPo
FZk0P0dMzcVETQKuejSxcERwEvbmNUiAE7S4D/sYjHSKo8dMTwpoffYOJxkAEiLYKw7GCyOMhWib
5jVEWqf7HA1uhVDqwEC+z2VRU9dAwc66dELrgz0WPquH+ikq0W167+aN8yEvAkbfI70N8k0BxLiq
3yJpQ3C9hr11ASPuETL4f+HeZJNCtTEC30kc3DuWIx9wHgc2FEhn8rJin0OdTu/epNj6X173euX4
gMb4P6B33v9Q9mGp1a9TLVNT/IdivnP7VbghpJsmtqjB4S95qvqaiA1LbyoX3eOzz08PWzlsMS+Y
0wr8u8KLCbNqSYIXbYoIKSEnnx5Se4+w8anilHGBUES2fx4fiKxleh/eGJLiAYV7GNucgk+olZEI
mAZ1qOuXwWCC7NzysZR0Y66nQk2OtzXdTY6z/BxKM8IUvAvECogbFzEzrGr6NnV0AedAbepOdt6p
GCIfkT6YlMTaAD5iY+uKXAz+X7D8mkuc53f0ZoX8/3OpfYotVmvSiQWaNSYwt8XEWYWZEUHy3eiC
R7mwcQPl7aKf/3GGpAIIjc29GQ6gIWoIy0opiTRrZaHkN+tPyOiQzeV9to3BVrAIZhS/B5FmdcP/
7qQQka7h4WciJ6QkPautctT3xO9TvadpvwjrNXzCJRBudQdCdncx9ZAY/UnQa1mxA4SokRhl/Jib
TvRTh8IG9A9vENqqwjKtSIE3cIkKPaV2ImjAy8YulBHPEFUWjSq9GtGtUeOV2dHATHlPeMbwkVvy
rjmGgPbV4VgLu+LrFSSHyM4+yNY8K/QJhbX4aZHz6wXj62Ykl1cf8N+o8iP4rqAZCR0AS1K51IK7
Sdgaf9ErxdgomCOS4gHCa+U9SVflK+eyNAdXkUpX/B1mOTKiDY7ojXq32aRtUv/u+aT7wQjZ33k/
nmCg7Xqg7XD5zfi7K4/rxvnR/HOxQIa7eiZimmBBa32Z7rTKL7ZvL8SBRZyfEzdTu2DrwkS9LlwP
cqdY+WSjJQNMF4RX1oyNcgYPdGUHdSC+gNdm8ATK20VCXJDQgIL0I5jhiPTfr9CV5JEHO8uurd9E
2x7RHSOaMIqTuit+qSgNOrl4UNYOxUCZKO2JZ9O1wN5H6WtCQUPYQhm+rIaGIQATc6ZCQf/h4O9B
7dG0iqYBYtd3G7fkMYVu2p1forBB/MxD9/fO0KujTcU327dzneCUJ8jVOB0trt90LX63V0BWtL6p
aghRMlqhl2NaSc1v1BSaX/7NfNmIOPBlXfxJ/vM7WwottGT9MLtBXVQDbLVfOi5pttuEzJV3k/RF
6U+RuRp+VUgpfFjbfHxdWfAk0z79/g5y+nhgc0wfNBxE0U3R3wCL26HpmKLjjiJuyZ6uKv3BsUse
gRvG34sILcZrPIWW5+3Nnkc3lFgr3sGlk7JSmoUf2DKLWcwaCqNKepTrG0iMDiOdzUaRhZN+/VeG
yZ1uv6AaNPzjhKX97IiJPBZKJy8lFzjORoTJGQUYAUy/rFuLlBFsf0pTbibPW/leYyQb1F+YkSVf
Akj2mnTKB0mwt7v3oTGa882tX+fjdqwyXMvNisrM9FMJmLbej34Pisz5YVNHWXPeKXp32zXt0/xU
YIiVTnUol1xZBchGd8eclYos74mfbM8CxOQ9QG6FzhSrlS+TbgqcfCjh98XmbQJ8pFlqEhxyq7ls
/AtGtwQTHle8EYAP0P5jw3IU02smVssmbxcvdXAJ+lOoZuVKLgKS/dE9YCOKn/PjxaeEv909H9qE
51VvusK9SLFb9rs8m7w9tSwxn0+47XTR0P4oy9pIBcCKcF8AUaxgEXVUk1fPtS1Pdao7IGWjcGQx
zDJbfe+ETTLakOVkbecmp1kLa8IuVYBlXKoT3q/lkp+71z4KRVBx0Vek85oiIIYj3mWhtG/PMEvD
mt0vETXRUoo2zDTrVRn7e3GQotlpnYJhH/XqyucsVpimFKupWXBfD7dwcBdc+3L+mq8X+0bwwZBZ
Mzb3D9vabCps9syFcrV+urUImY3i1II1NGwRV2CMuryMIqw1SnGQp+9tyH8yatlNr4FFAfFNRjiI
BQZa5q0B6RGVk7Nk8MzLh6++bp3rl7wdnbiZWVZ2ftZmfKhofgkGKunaldQsRsxx8XQ308LhkaX+
fjgLG5MJj21xk4fXjy+p5F/lJuD6h2Xr+auim0DWtXYjfaamEN0rMdy7vVYAvKlparrVev+JhUgN
yJD8VvZNUK7fdZJR9bjhA74JoPansM5TDbr7FBBLFbKRkIsJRnoc4M/wdftUkIbiaFRCc4dRmfQb
KctzCKhZzBFZIMOGcF2gBfzxH0qPzImTi0nJW+7JhuUYTL6QHXA2dfVH2QzuHEJOBp1L8kxVJ/J7
6ZcPmBQZfimb+Nzax9CgAlTQZ7AAdJfk7kDfkesz1Qv5C11cKiHdS7fVpaSK6thAbs1uqDNuEWUj
baXspUnK6f51bvSMXzsE2VzLUyKzJPGVXLxavpWjhd3sgAzIPkkzGiZwfPWRQcOATn1cE8CQE3zh
5iWJHAbQGsbjKA7vYeb4XhkFWMJW8BLdWtmTyA5TgKD4DJy6lpJi1NF5e6ujDspTUeFBkfTwmRSG
TKW3d0cykl670YyoS4bQQiB71wLeg23WxQaIOmfHMx+FnQfo4L3kweCD78+zomV9XKWzTSRJQXkh
Ad++MzHy592kASERCYclLn3IRbW7jWzPDg3Zthh0NIHMI/g8l5cJj99Qk/elFf66QGy6ts4an/dU
KuRk+rbwTiDiBnuiXu8nbtSONB9t81I0OvJ/jqr2gm/MUJeHLD3zEURAZIGZAGQ5gTvAmHN8hx0z
3Ot4n4ArrhHPfh0/a/nMj8YGRA44XC8V1S2HyOL/HWGCk+TPYhAXlZuMz6guPZ+nCpSii3DWj8nS
Z862agD/hNhpu8kGHlbr80QDaNFzuyFiKj54nkese5C9nzaxxRKhjt9zUFL18OsxJe/5RIA1jnIJ
baxeQNlm8PBm8rjxMAdamlya/26Zs3mviEgwZkYvXb/lBgAU7cJT4vQrFzVazZLnnkraIV4UMln8
bJ+jxv+W0QOksx9z6wI1jEhMfyAxaTlx6BUcWhmqpYcu0wkDVQL3pXW39yLRXniHWhJh+qqQUwM+
TpUAarUBHTF07f/P6m6T+cXG3GJYBBgFE6/031NgfnshGGAvBkrFOZ4+IOst+3ZYyHaeLRLaDjoi
eC5nmFfhh7Jcue2Y5rSsAVcxSH1E333G0i/KP+k6k+JuzlKDHSuCgqUerW03EHEjTEYMgcrNXcvy
z3xs4Dqq7XKOBphDp1JSZ2GNZUgRUtBHnts99UhHeL47GvaFGRU1EX0A/0LFxbXrq1ir0hMbH1UH
z9JPXWxMZMn8A3qgyEE2alMRVIj/DAQV6ZaBvsYYjIVtvBOtzBlD2u82HzQebWrRC3LpafChcYhv
42WJ3TKTiNPFoYIaUPfmCODdhiaarWS/zLDpgx7c2mY3wKvw6khHXvV0/2HC59cYgdPwpUinm0AE
r+L3LO2ZDFMfBbMEAlnHc47PKUj2WW3agOWUA4ZzcqzF52FM9TFTrFKmwLyCKTC9huKpo0tmOds6
xkVGEV0/QA0KnvpT+9m5IQi24qKOhdye5LkpnlUlRDFeAxwMV91iVtnPl3l+hj7cF3Omk6vkMr9n
u3bNwD4uZaKQSnMqInRy9/jSdE39itGRT2wnGyCiUFA6kkSQoKOw8TvkXndoT1RP0yuDWK6PEhaF
MgYC9DzbIUBcVlPPKSUlYSrfzZK+C/BrQgQA1HPMqfi9FZx6FZAP5NvlEjflrcFenttJBi/T5S/O
KOvLbJEmFiuX/3UQH5oeUbKQcLNwl2l09jMUsw5bu1Q60mLE45pJ1AuJfx9oEzvO2zpCZBJkOosU
CcRn3eaYB4qgmdoDG2LyQ33MFF4BgEwud7Hx8QoqkzqJR3z5uiGkpVH+pdDWjSu5s+hWgRxRr0Un
MGOjNGZUu0Txy/XYQnMy6ISViaFDXWaoL+bmiTG0PI5a2UjP/TvwJOJIif/I+MLWnV5B4CHwRmZG
bNu+Snlza0D19WCGdWN+Vb5Fas5ga+ODswR/CFmu33IU31K+JCKai4QecPTy+5qCP0ZXYFzqq4xs
XJqVZcunKw2jgPEBXT2XA73KLApEzKqnhzSTX9mTPQKPfMqloB9llFt5AO+ZLJrVySl7RGu9qAok
ukUg7e49YbX+KFWgTvOgWnzgk5XhtUijzO2FoJDKHGoDigynJWzad0QDMPs3gchKiKWxQ4qDarGM
2JOG/Rtv/Mj4EonzgVrFdSDJF+RgS5sIdNAt828ie0AeJEbVswmUBULOpD6xYbnZUsTgX3WfD348
2/kKhA2MobwnoD+0hVyXnzGEV6RqNdTjdcIAZLko2hqlQj0ajNvVAd5SrEBkuUsvp/8QMAwK+iLe
yw5f/a1JwYZVrpvsmTDlhxPFH5e89W2T/TBUNyhUeAOu4FFUiKNb5q+WYotLoRf1HPy8aBe32xJN
d+22XkkrXilpYHzVVP1LSWQSOwrG1B2Ns/THKTxV0scXy4mNrCErouw7iO+gSFSkFfGbOJ1QzHoM
HqZa3JJp814ty76e8bJFw1diVXnJZz6wjxbt4kVj+AVA/RWPaeb44vMLhf6n6ZL9sB7QMj7/MQUR
CvvMhvlYgbeQWhnMXFbMFxGe/kCWsNR03WBObXF2ZJ2NH5CFBa3EaO/4hCDfl/hcVOkFI9RkUdMt
ss6sdy0Y+pRVyRAaJ02c5r4w28r+HhWtB7Bo0TxVUxUauEz4STd+anz6bLKvv0Bkp+rxLkswTkDT
ejXaxxPQ4QJDq/mry7dJHRKcvsUl6yImbPmxJeEbp4Z7GWol4GAKN9DLtf8IQ3iBVp8UvSUAxXW5
N/HQ6GY+ZUkjg+y1V5QgtaLbJEyoFX/btrg/rIVGU1ECKhZU6TkhRR0DV3dBMsHisvm9pHcTH/hR
Gl0l5mcCEvOlDmB+cdAqjgZOfDN4eAh3CqMEbtspK5eiZEoKrap5jeYwcqV43JS8zF+rDshpl4LR
9jG3XhUWobWCJxBlonPPwmHYjf2Hu8MbVduh1auHtdpPxQJYiCP4IhiFlhAaBnNorJ2vQWMMNPTL
JPo1WKHqMatsyWwvfcmr+aeR2c3JAvZSKmgdg86rCrC2OYjwGUJZrOcIU8EYLmLlPzR03rNpV1k7
ZB3AoOcSwjsP1IDciVMSiREHxE/DyKJSuGkbHxydbkpVO0+Lz9rzCrXJ3faDaiq5BNtKvuxDmhzv
jsYMlDEmhk4U/66YJuBmtURi8S3ArxeL4V1E351OraoJBwoIQ7NieVLhGBWpEnE+vM0vWQsstX26
lcCpeEDDh4gagSMLa9kqNmMbmY/zmmmqMJ2P7RlnS0P2KB4sHlzrdXxSRbCRpoh2nL8HT5xNlDaL
PmWKtEbY4eGs+UKqfB1OlRyK8vSqXDHBkvOm7WsSck0aSB95Rh5MdtPJX7OXpA+q4rQl0Rvz+1pW
wT1gQ85i2eREKe9Q61kA4AU5zWT/BG3TQV7Pf/Nke/3WR7PuH1YGC0oq/MhnSOHtRio95WXmrFAx
j8KKtKB19LO0L2OAtN35OIYqil1Sq2ty1cYbJBCjFx2K9aCDSfDV6PIRQC1pv5SaYGHLYWOyuD5c
swr+q9ftmv9YfXeMcJDdv2B6E82daTxpFe/tjWlp/mMQCzXW/Qb1PaLmqv+oPpES/VFOHiidAoSZ
BkCpp/aDuGb5LIosLw8oar8tM9OqM+N3sjtqujRBAnlJl6XnpYFDAxv0zyXFXiKPrc6MFM5PTiL+
JTgUB/oBykGbFshKStpK9QKrwSsU4+rgleeo36EqRJjB5HPkFgF1MStwjPumHQlRk5tTGoCczp2k
N8EG2kNeMBuxd79mFJSONIxP+R2l3jzcgVxfTxpPg6UcwvH+LG0mmAQ2dVOsteJ9nVg5Vh3tzANe
THVEhtFuJo2+4LloCv09sTQ9q37snjjJa6j01VWvIj31rRMOAJ+dnQTlz5IlnHRZHmhB0KrQBQ6d
4j6EIhUAbzsSW5RJSUC/+RXypjysF6R8hHTFHz9Vbxw4OSrFH9AxL+Gwwk0LrUCq0LLOiHdHQSrU
UlBJqu99rdMjg2sVDZtba1PWVocAS4oAGE8IpceqbwIXD7h4dCAglTiY2dBrwwjjSc83pvcux0TF
WkNkL2ZditBkoRJ6SGlgxc+mpWzwOQfVSHJIShSivaGIFHGemPGvFeSqb838QcwPK5nrvEBhAL8T
vu34RdM7THd0d8UM/ZdQdplwPQDeBUkN1mc28YSm8AuwGTh8V4u4G4ul6NUUyW/p9iMvs2b5GlB+
UYAEPqD47EnKJoCm+NhZabqcfKktlUKAVK/yD9ZO7sOfp3+2m78e72jU3AvT21mKnm+aN1BtgQnJ
qsXhBoUpDIcWghjxtzAs94OXIC9KZ4XHaBLMvfmVTPdqfPRXXRN0NWCrWuRb3MVtrxnn93MzbPeh
ZJRGUmm5LhIRQQfj5btd9b8KRR8JO8whEmfpdoPCWFkLqcXPfWxtsWT1gpWWuwJyAVP+VkKLLTH9
PXMzv3bqOeP7ZTrTsqqAxnTZejPpewXJYTl4iGRGqOgIwtenDXeEcU4P9HBC90BLytPK+/yHU+in
NWrZCXawsW42dCl9qnnp7aELdatSyzz+DNlfbp7g61KzGaGWdV7QS/DuDzQ1LMClUeYS2FE+caUx
MGJ9GWK+Jj6rJH07IPu/zrA/bJxQNgIlaAuDUROhRrq6Ru50MACZj9zgtmNvjbYEJ2jQGgF5KGBx
uwRC+Ks0LtndB2GCuUmOBkLR/SetxcMFlNSyWb+Ym7V4kMa7Y0T+xFCr9D9BAsR9LjKnwBGFY9iM
ahtMK6nrg+QL3ycyWe7fZ44CIA9MsmPG4TSnNS0Z+PV0aj/1R9UbVUNzgnQu1754FOy7VEFwST45
G7KT77l8XWX+8TVM667117hxsx00GC+UPeKY1zG+G+s6rnLbCpmjEGzo0MKLsh7sIOA23BcxJItO
3+Ar75s5CKY3UvYYkCGFecQCl+WgH4J++d7h8ndDmCsJr2QgYHniqun1hy6uWebAfEpr086D9nbS
Zy3Oy+3v7XRdW9yQi3csxP7+Ss7oHlmFm5zIjh2SmscaTLqqJuMPLIhwHUIeyVwzMMNgqMOuDeS5
UeeDZLt9kt4VaaPRTm6bkeGcJv2BR2MovThw8AfJf4pSUWAyQjwyj51MOX+UA/VzSbDwPFubbar/
JcT78dYXT7NRZR7HcDC1ZZAWirY1N4NZVDsQFbJzxvW5VGPUlqPlVo8GuEj4W6FZ7m1uEb3LnAq8
iCL9sNYS9PW1zJVdu4QCd3m4NSp99bg6L/QFhv5ou4hi1UZnvOPEabLTHFvu3p0a1N5g94b19trv
FMlRMGFEd1UNnarYk8c+mtDq+gZmgO3Ll4Qj0ZZKbUlQJZmMhfnUKTS83HHD70JE0+mCT/BIssE5
AXIYNZcEJQIAhboczzu9XzCzTiHQbc+ONhja8NzZn/bl4DuhEoUPc8d3ZlHuMsuZergrLbOBuyHD
4OaB4wKpqxTz3uQqrVjJpHePYByG5D22mhy7XIOUPAALUCoWrXfGl1d79dBiNnFZQ4z/ZgpRAUjm
yqEW9lfPZyY19EeSU+kA3pR1vvM7bOXpRGxbhgMISmVRibC0IBYXzItxKBdOtqaBZS+XKSGiyLb0
99KA9Xo2zG2KFWnEeAl5BFSpqmGl6x6L6XT2QKJbBtPdBg4Yc7uIWNQx0XWZGj6v9DpfOmk/olRu
UzRgw31wr+3jaHp8zASLEtLvgcnDbKkLDl1dK0e933Yvvulzm3s+ue8vcaQTlIZV5rMVXGmd6USQ
71IxEstygzApD97rEw8t8ZrEj/s24zDpYagH4l6mPEvi3c48YWsXsniDG+7QkwcgtU6Kx/J551cT
DOxzv87N4+yoKOtF3advn0H9EJMmJiU3Y61zcjqKsoYDCeiGYaOe1z+9x213DbwvywPbzYqwe/cU
ysqYVky4g9Vo3sIA6NAbepuIml1J3F1cv9l95yjDnPQMVCEZ3co5KyV/V0bi5HN2Bcxg4gRwnf4S
RT6ymfILQcpaE4ebop2cACNah7nQ1dm3tVaOsEHLGbkbzgZcPiDxdw5zoFGVqQtDHPqB3I1ZrcXw
PcYprJVscro/FBVPPtQYP3Sn8AXD7lf9fZQeki72ln3PQQAjDqYBzNL/1O3NoSPcAtYpyV2/pSnL
EmrHhYBusum+FOSWT0Gw2RIcv2Gj8azxiSrJieCOeHAKD96BDzM4S0DakYqipee2eIPuoj+EYzMK
+4Do4PJK4JTaenB5GYMng56EVtNkGKFf32Z6AGotW38njPyxP+kGafWY3dQOC5EffKnKBZkMbfAB
T91ucTPGMgP+PwhzOp66YkGM62M4rn/lHy+6fSdqPGsKzxRbrbyp8I5juJmFkm6EmnYJyAFe16V0
fuSsYyQqCZbZyD8CQZafxw2Ia5n1mYsGzajtpfekBk/NH4lmiFmo/uxG2U72JJABZh7VzmF3Msq8
r5jqFv9kdLWztFpNgTlkLzDm7qiP1ljPJoJUWpznmmtWHfNPwO+XRa+/AuVUD5LqxVzS41NthLLV
lmKr0cLhfV3UXfo+L3dVouDQeoglpDDlRbCKgphe1JsN3Zw0+7DjfFSDtpy0NSNkpufnF5zYXMp9
2d+/f45Yhx7I/wTuefZFTfDYiE+LGYtxUNpHJOx5unTptClMLwAPC1PYqR/cmngCh4YFt0i0Dk2W
ZefCMq6hN/D9yLaFQu7KQiHOAb0/5UvQjR1/K8MSnQ4XhJlifCOolXrK/htXRDJ2JXS60Vl/tYBm
x/OHsLmbepSxriRvQ3YuAULLwoK7aEmrlPBp+OLm92uLqrGI6WWLKoHljFqNmAwAdSNqW1gvPaA2
GuzXn/lLhiI+DlV3bwtUhyo1YCygSS5OxH8M24cuKW24ma0pISBXHmhCmLUsnRuj3zAm0/p2zQCa
3BnY4L8JdXtyvPN9gU+cp3pEbqCKXMbnontLTebi000foUj0+tYHfKB05NLKOC3xcd9Swd7EtZ8H
VE/XjIHHZ8I+Ne9YYmZCew33ppoQOCfKM0c7WQdSBn7phFfzSZcAHhFZUhmrPeKW4AwXuJQUxm85
Rv5XlE2Dh6CL+ezJIei9dorfaKKuAK+qiOvxfT6lUoD33bgqmykRrwvDiq4EWbb7LjEziYF/09tp
rccdR7W7mvEtUtoW3sRPpSww/Way3/bGRH1UjcAlCtFWck6Eum3MNH5sW4S5JI4mL8kAhAinl9WZ
Sd280RsxlPcIjZEvg+EfuHL00NPVBsYW6cBd1U5t5u9ODCx4+9RFf3O2kxXVAOqIRFkHY33QUOWE
Cn55fslpOwgTsXXM3tH4NrygqtxrCVEDlb11Qe6Gd1wgHOi2qM0ZmaFMYOlHjv2CggP0u8lbu0Q6
QGhKqOBfjJiHPuj3EQWVuMvaAyLM2JHLVIaQ3fCejoLRjp0kBOSjTvkK0rXk0GLXHkTgmm3sU9v2
wEWjwsKIik8JK/7gdnzjcWDvYDrHfZlgIId7+pScsxF3ywG/W+mloGAkC9nj7I1RIGRf+Q/mtl4Q
N317fhriod+nC7vrc44ojmF+gzMI96xZmg4rLdq1E76l83OQ9pXBAEsRO3OmX1mT6MrbS60KLK1c
jAhQgE8G6yoGTf1Z8c1lUGQ6+awPu0tARySGY6G13aBtHkykboSQdQosF04hRWK7rd+6U25I3rlS
DsLNkH1KjFE2fLkCiqcEwcnuwuGbPxnowNlWr13jYkaTr4tb8OswBDQH3+RP28EOWHtIeL7ORwfx
kLT+VhUEYRdTdt71BD6nxB1L8YWEQFGBdrWTS0YcENulCeaEcEwhWzMz8qyFrGQTZ/UNGTKNvOHw
+fYeXyhR36Mk13HBQvCsy511VAKzf1I17qbTW1rI5uoLC3R+3Mzx7ZfFyXETjDqDBBh7Y1LGMlZg
nUPY62aW5g/IltFXNR5DkWIwrxwugLm/m2dIpMnbVNelw//iFdh3m865VGl8zGUOmxb7fbIee5Sx
Zr9n+bPspVp+1pNEJ9Rd1vaa+5CP/b1e5j1vmS6qgwt8NwOY/tzsf7v9CAn3+B47ixc8NxiRiI9G
KVhQKIOm5eNwyFYmxGDUNx8fSibOK3f0ccEGsc8BOV97EP+e5+Il8UwpAUBZ1/sNkW3DNBC6OUOR
OX+9mr0psO7ejOhcF440BiE1OfhKKXMHpi4inlBzZ1brH0ZdeUXRII0100q2KonCG4MrF6Ga4D25
iqf5dTgnlnNK87hkY69ghw3E6vmJOQFjUshuVFLF4/V2SpyMzdOrFPHCL7QebLH40qRYw02QevrB
+umpDNt1YqSF3luxvHSeligAQbeiIqgpGXe3oNTH17kHpbGF4wYlEdQ4+yQ1lpoynoIm/TQ+tjD7
AdBmWRseHx9nMPdM1GWp0pIVWZnGLOOul6uEYLVBMm/w7JMqf7VCytIhneOYgAEHQpfX39z+L8+y
obdSZE6xRaQaK29YR44HEZKjiMzwf7+0vyNloPyLrwAdTm/DxVuXbXv4U3YeEtebb+JYsJb0bfKV
nqTI9gcPxKIVpxtNEkUi6lsB1N57Ya49GYAoL04+wVhdhy6ePJk0+aDJcnY6J5e9P+BW+91Ht3fB
pzr3y7JvZCuoqNTFShgTa7tdzCW9eUMaL/UTa4fB+VuN5s5t1uMvBxZHKmdEifpUG3PUJuHqIOXV
CtzS3jBcoTQspUaQZFIKsq0EHIvzXALWpTbCEvIA/Rtv3YWn+PtRU3rr9s+HiCJfAWiUyGsUFjFM
Y0vSQmM2El2XHi9ddxIyO5uw4gPU0Zl1punRx7rhL91ONVjkimWh/rSaxVPt39HPItnDo6SRWkzo
26/97asPrTyZQewXvEAhEgvzww98BxZ3IJkziiVAOd7RKg52BbJ3sL3WC+VsJ0msVhgDdEK48Ubg
Ye9ptxtLHDtLrgjdNjFMrEXrKxVIz0Ta7vFKz/M4L9wIeNKznQwpqM8AIhq9HbPNQB1x+SdsGRLj
WbsOvF3AHowq6pzRrwHUG1FVkMssVgLA2GfoTBbbS0Ak0wC+jreP/TG2II0OE9KjLdHHhvAOCv60
wClCRT79X3HKJemNlr4SRd3KOrOl0nNGYnB/gyuDSDcs+lVbhIqAm2jZ2KzXiBPrj5K36sKDrgjt
D/jFuK5KTydG9GynuExFHuirhVJWrbLzc8Sjs1iIaTrBsJc3OdZ79yby3f/RTgvnMG19dMq8VOsZ
d4Eo2NO/SicDjQ9XV9gRwicfYvs1q8InyBXO0blaAKMYQSw+OlvN67Dk04g+SHLCE1TbWta82k3w
fKarky0jNRHm/MgjlMkE76X6Tkbm8YIIv7CvLlq3sOL91ThdHOzN7ZOwjFrrsGLaGGr+wYcVpHs8
JzJ2Yk8HZN6tUSF/vAHNfYn/0TjmNViVV0q6ichDG8w1UDkjQb7vRJj8uL8pXvnNGRT9bChlorI2
UqGmxVURUUqGY6bFOf1o4aFTbeF5XPeQh36kIqVfMCEPnmIW9Cc89G2b+yYG5+I0AuekIhHrZu6W
/uNvZSAnOJCtZMXCRBZeu7wF3JTZgdPGDiJlQaJp7/QgvUQcxQI1iOUyiPr3sfoQttJhb+uk3sDZ
X08g4uiOfMMeIc8HArNJ3KcmvLivwsFvKdgUCtMVIsTbIrNrTXUJ51G3y/pjQMzUj9uf6Dy//kg7
VSOAfz+KyFaP69+dH8wqhYkEIBH2SstLx5tQlQ1WPX0jh4a0JZJKpnjUyTdqokm85YG7Y0XeroH+
YkdGh0troFTEydyCvQvkb8tpjshpz6PVDJhTvbGi09n5grLSN8TgFvvqHX///i2upYxKlDQq7nRM
VXhHsA5y4XdoS4LFTo/xumtXdB4UTjnqB25U+TDI/GkUDi0Seb0sEuUb4rCI+MUvI97lfXxGhrM2
CqUCQrZ/4RbWLEeCJ5LLcDDfrsHeS2Z7skTk87pHVyzCxBhtH7gH7RbjVE93NSd7wx6vaNBoUKZv
XDqbQ6A41mZhNrEJomAKXWCbkpi7hB3FHmcQl7wv3eMbpP2JsH0vQ8Iwakve2++du/bUTZtNJxra
6teX24B09SPmHCL9FUm1Z0s67NMtBHd3kDVOvlZuqov0hLiMoLWq+6Z8Xf4tegzWeMco0ZSaDqy/
hFlDfLOk67ImMtaRlBrhn8qeV+hnuS3kNXDDeD8fsUTwIfdTqLzObzWRtDA1ARjJt9ZBi0abLPyO
aNPCCitu4NvJRdtXvLaRBQhGVtXyLxAdQLRYkZy0w7HWlsbSasFkThiEy8zqPBE8MNlTHyRNHXka
3mkt+GON0fgSeWAHI0QbEcJuAqBZtITxn49p2671/9E5VU8PAUVW4mmDlyKnUEUJyuMCL5KKs4Zc
WcMvqP5nC0eLBsMTDdAQnbS8L/P1Wst9rsbTT2DsKntniWEQI45oVEhqNoXevcNabCOxcrN/3QdU
CXRfIYBFVQ0rog/UwWLkW7ljregzo0iDIQVHqHNmQd5FZ3lPp9r7vYKPvILmJEuuo9PWINxpEge6
N/HY98s3ali+0+rbt/Xutj2NPdIM+kyMq+E2tMDZTFQYm71hVky63JFNZ588SkHxEHj2qqH4EHxs
w0FJ4+lp8w18BivvMi2WbV/bsba72hCCVHoiwyENNpqxmI3iTQIPc2wga9cb7RwfFdYp7IXU4Fih
zhJOcxPD9QYdmrqRYHnO+YxjZ1t7T/M0X4G0pkJOogw03TlJm3rRG7q8AeVMARwG0aLy+MWikdmq
GX3mGsLJX4KpLilpq1GdhRe/DobV3UJlNmsuw16S/MEb2O+wK4UG5hWzpxVkkZl/qNG/uCOUjNDg
RRKvYVq9tgP9vfLbEswboaSgY23W5ta8nR58uWoGsHpfVj/45W7NXEAWvzQKn4+G0T//G+GGIo+e
HlYHMXJpZWjUAFWBu50QdCICbry6mIyDlEu3A8AV61X3Sat+3LmMRbz8Nm3oOmzZGC46ngSr2gVP
wR5IH97RSGxIbAdQ1YcUzxS36FlK3BJGfHkgUma07fCmflYUiLgJOoZzOrWIizslqxuOhjHMeTNL
ZO8ErLqjUSsWIgzsokDh9NuLsyeamAxdOaloWnufjCqqYv3WnOQTezbdtsGWezyRJ1lV/Sty0bxw
XyxPRjjWkaz7nGBy2+siHWyATqQsaYzQ5ELsbfZI5PA8fdB14NP+T1qvRSoNcvQ3vmYWBT6ibPBS
C4sevFl9rG9oi0nJ2d3hvQeq6PrlQiQ04NFqEv0zxfKPsO3mLQbhF2h+34ge3I7cKGrxJryVHi98
9c9tgHDf/+tCJBmH4nfaBrVZX3ceIeFE0uBt62CDtrHONGuYiYJ3eyZhcEFgfCI368uiWLOrFokO
mA59BzI+9TtHOQe04TRgMdowORle81Kl2UtUU08xRX15Znxjqiv6R722KN6XsvDVMPqPhIWoO/iK
x9GClsSa2lryC7GEXeIY/h10E/IU5T8xSypET+zoz9IZEdjasFT8xXbiQzYMWpoaONYI8/B9C6/S
tcQa/Mrnm1rPaq4mZ4tBXbveLrwmchXYEeY2SBU1dhhcKoPNErGYHY14USdb5dx7iP2dHk+x3xVB
WM5BxB5MPSZLEqwh1X+8N9YPJUlS/fWAPc6GeI8jihnYf1NgOHGKMaf3F8BZhJEPbDYkw1M0Lpo+
zs86cfrVrOL9R3tR21dS4s+4f+/mRSZS9Vw/0NdjXjpzjEOdgti5V70XPFSIYjt1hgThgtk2/TyX
sxbebJBR/26fsY9SfVd5nAUW1k4B0q68UbwOEuif/nEgnNjlnEZbiU0hW8HFdy1wNKlGK0rbecHw
Gv/KwYuDhsnaVdr+nWCZxdxrz0CB5+mhArltqRE2oc92tyyj4AzQDLGFmChtdTZhslxiNeoYzsTt
8HCW1X7hAUEP/8GtBs7IMhBGXj+xKq+N55RpilIe3ALXodikvE6Nl9y14WkztKfoMGGxZ7ps7V2q
KCvepeeasqTnACmTuDhclTvbNE9zBGnwX+rE1k+T73k6ymhgwgw3WtrP9F012ZvUava+esn+EU/V
BE9OxWcmVgE/ac/+asVJClFXuIeBg4O1V7Vm86X+K/fiLl4D2SeZNtcbLSFDHqIz9j3feBl6nckC
B3FbdUsZyWHtYucOtLde00oZJNOkhehN2Mr4clD7t8MIzrVRxoIDw4a1JvEn91usFb8leqNg+as3
IQTEx29rL2hW7aYlI+MDuPERg/DBQRZ1mPzhu/g06NmnTiFW1RzJb3oHcX/o9ADSA3hKlu4pT62S
lUfsCO40GWs0mjOhY8UW1ftCQ28vmjhyeuCEKIGx0BvzGc8/YLXD0VI8C2/FsXG6H+su90h2U8Qr
z2vaIfbHnZrOrBdox1X8HaRsyyttVvoyY1KqXcBmtza6GZzNQGmT7Zs9uELUaycvEAtmpL0vwEx5
Zf5LBbKRrxdkXBuWhCAs2m+YvoAUG2QnsDP4t6UQmZ4+TGkdJpRxJXLyC/rm2rc177gIBc4X3ead
yuQz9MW0anvbqhDSu0o3s3WubUqngai1j+jlUlUb8b6vzHl6Ce5peiuIgtxiCFBMKPCsJujLKDwq
ZyxGPv5Toowjkev8xh3B8XS88tZf5udIYXdJJ4HIHnqdq8R4HKdbuC0HUpAPCh29U7YmiiaHDqx6
7xgjQtUfpEgOrKX6rBxK8BO/4pkuDNWxKvGKniI8b4ssobbNrc/0GCJqZla4z2fNLlbMuN66GtJG
5K34r9PztmkgewOFvTW9/K7ylQdVPUjIpvLHiXjd4H9KPpK9ZSFvM8IAKWxYIIfySQcMnwpNRK84
aidrDjrjXejzZL/8OW604lzt8MmiJS7AkKpdfkBX0in5/PJ+SvnBZL0lGnIguNbLkDxG7OgloKwZ
rywyGL6XCL4/2GAA5KGAMRr9hxrB0EXauAFDYjwBFNVK2xeKjmTXKfjxwrQZSei1nz1NlfJ838ZX
Ha0HffdddaxCkjebYZK+UikaRXeNTIj2oRKBCrombmtCGcvVaSeCsuVabLE7yyiqZHctsakTHYY0
nbqYLx3/rvNKbD7hCdLajo7gBJHGXBhSOurI/SURlnoU0je5T/nzMx6IqlOlOffbE8YXVQJfs7WW
E8Jd9P4aIr0eMAfrRqvHU7p9aZea1FR03XbECDYL4c0CaKCxWajAzotpBrv+HM8CHpooHbk7xNPh
82O2K3skMtI4EL8jNNnPfYe/OuF1NeNe6fZDZr2nKbKqSNL04E1OFH82CK4FLRREuxRpCJlBBwxZ
8lJj2hK6lr2e0lW5dFbFj6sRbBcjVkiLqvQZmRWLZMIkeixfIp3IG+7sdS735v3sTZ3goBomv5wW
IsGri2jcRKzBIdCQumpY0qPztBKTlPYXofEfk5YJHG9zMphT6VkpN2vdBhiH1Oz54e3Ixaakyw8q
wIlwjnt00ch3XO9nurhOlNtnpwGoz79QrAiNxT3XjwYevutNIi1v00VKiAaP3pzhJ0LBBeleBC5U
rE1Cs5d4MinhkG3A+ETti9mnhKtm9XFGCOjmgYKNjT/lW0YMEP8hB3lwScqCePTNQxRiyB98zV27
X478CLkImPniSeE6WzUoIYW2j94Mi4O9klIBJRowoSclXnC1wxacFvRnHvWrdipt6c4qujdv9E49
Lyp0BoTSqiAWBFR7dlGi2tZD4RdAMvgQtQ8NyUUcxetXD/SfSQ1E/WPR5+9L7tGV65sPoj6V0Ixd
stPVLrUU8t11QLaJ/2wE2PiT/qHgpYjpjtQ988lglX7AuD3RfzC4MYW1uQHwgms0fuE5v3sWnfvA
OYR+o+O+eP6/wpulaGAyr93my6rgIPFvOKoUYs24rPNQOnm+C6PrEb2amDDS5DuGPELgzb2iCNMz
BAcyzwF/r8fwJqbdObfMRpQtiqGrfaK1X5T6/UUqEQdoPm7YOjv7JpcMKOseDfB/rYIBiYzo75gw
X0nX+zZ6APZecfunT/Bw06pSuiAeBMwtvVSNr+cV43gLVxK0u67E1LQ+KT/8rivmGV/wqYPa4VtG
FvHShrTHBkomwei1OiGhJ1HfWmstcZtzRyXYx+e8WyWjKZAwf4j+CgAp+kJa3e5LNeV8fbu92/4o
7jCwW2HeHQ9nx19vy86blp7BLn6PNWfDmQtcPZGgAkioeT8cnvX9p0FwAGyxC/sag6hRqIbk9qCH
KXjIBecwZjCtKwaFY/aRgfvD3BLuiz6SSeXLPwPXWcSto7l7G7h3rYin1b041i5FMoAPIHcc5SzI
zW9bscgyFDa7hgvZBGRKIJcDS/h/S6oEAUx27YdSce5PWdWlUAgMx11dBQDkgqTmAyF++EXfx18E
udBtMokZ/PJVPTcS7mqKpnPOkXMio+XCjo3dkyPgHoaOuAxMZ92ivclbaXwEJA0StFpxu8gBtGMO
1EQZ+G5znTdN/YspeM5lqdBu0UEQFuBdfH5HfiOClPlg9JObG8irbkljFG0mWnoAwwwlJxqWgiGW
rescBOzHvFxKYdW6+2sNGetx2blX+3P/2WTaWkVrDT50NSHiH2/cwR7ORy7nNW/YtPcyxqMUGlIg
BNvlPZH147AZ/k3c2uhHvehEAPjZjamaSDM2ZnB3vgL86ALk2BkOgcIgkawl9UpvLf3Ij2MaT0Fn
7MJnaooAMp17bQ4ou00SJ31OUFlvOjPTHmxJKsAlu/ygbFj+IwLDg9CdtB2+H8DBAhkGwJoCatD1
+UO4H9hhJ9o6oQwUovubu1ALNUK+k1SzrU4I19cxTHvy1WQ2bD3OoIsK0dYEYV2B49+cHTr2R7vV
8J+vuDHEeyVvYrGJ4n3/awV/8ulY7ZHqeb0H5p+0pEyg5nsCpNokxJ1HsYdv2XyeK6nvHc3EQspB
+il5Xv/jW4ew4WL6D6RXBkvGyXNkPnhVhN38fqEj57mUmHL0XD/DWXNtZaITSiAWmZ0VkXGiOpIJ
zcYmYH+g3KRE93QVnaSTXmkbVhwa0n5p+Je/ZHWvN1uqdgunw1qI+hsot/cGysjuqTQYAJSnLVJ8
k7UhHC6LHml6pFZvA8tHDj2asK0iJ38tygREY3drXcLvZ1Wk3r7HG+/K15gWJtJCbeJN8CB3zYkB
RFwuRj5C6+6ZQKxT9Ud3IW9U1QD6ksrPCAO8XmaDvT+Qsx0hkh+uVXRSzf8D5v5Ds50DHbyF6VIR
AFcI7G5U6KX8fa2ukzVs3FWv3MBhZjZnjppGSI91ZgyQcoozs5ayLwahTPjLkWt7xXgPUqflHkLs
/JvYvtOdDj2pkTiANTpuK2hQzrxPM1iHcAIzKLuMiW/WGj2QOvkbwrR+V8jmaEkI0VFAt9PCYN1u
foWjwjco4Xo4hLBjDROpHsHfkjzV+s81AOg8pKxOlF8mdvaLdZr+phnJy4XduTXXZFxUDmFoof4d
DlS7gjAlzW9LRydbOMClZ6fH/hdZO4MsueSfC6g+QoBzDBvRg1oxincHSRXsuTmQLOlnLCe5G4Xw
0hRdTzo9kGHGEqEpZgZ1M/ezswkeSr4yGWHz9p/f9MxTgOaJZP7o2EIh6LMLXqtVpI4Q6McTNcqd
grG0Ft8nKBJXu70+GrHNubtjSa5bRwptfkssw+mh7N9OKryPJgRUn4kgfUk1Cf+7hjVnn/QPciGz
r2kjl3a6X+/ul5To8FCBP0j9CqG7mMBiGdeOxYxN56nWcvpSuU4aGlTTj2qzmgD+bbPqjKsxmLQn
4K1muLsJi6kwsgSOUIvXHpqWGrqcmTM8EGQMv3Zxx5U+asXjcyOVK4FsG3DXCyZXVkYeC43WuwxK
jOcTeWW+az1dizokByhEqeAAqF+pd0/TcTyZFzOXy6jR1sOXmdK949/3UT6xrwtd3ALMGqq/V+ra
+WaiQvchLoKvjmpwzlZi5y67vccjrZY1PhzBlhXf2SfXi1vZKOKwCFCjWxBiSuYQb6/ULBCTMxWO
An1fGXui8ugiH5ZC/DJG7byF5Q0FKvafY81UvoXe4aVb5/1LUAEr9w/kynk7fQTTKuOMPfdcYTQJ
V9oz872rNdZByzGMVsCzbS0VEoKGdvg7LfVbdywPT4/RJZYeXXx2hBVeUNL1pfTxM3XwB+Hgar8E
+0WuiC317Sx1T6JXOrB2GkYzfJGF/8TLODcD6KfQn1bC697ObrL4wrjHEZMLCC71XAWYWSnBFHlC
p/ly9MS/hn4DinjQ6FfCyviiPO2lbj8Hlu1cekmbhDC4ZQKlFZxPuFcTLeHFVPgrO3YoNn81a9Im
XyxCLF6K80k88v4+Vmwy1bNDf8SlHSzowZ9w7uBdORkHgx6icdMYVyEVCtjc3H/bC553PaiQLEsK
0zZpo5Ko6jxYMay4ruNUNZ+GBmj3p9l5/CV80SxNMoT1XWfS0FjKoAkJBVHWi4pQOrCA0I8xG85P
b+EcG5ayRhJ/wxg6UpEiJDwo6c0yKf5XZvGlyV+p9HxntHki3Qu7hToG5b7KZLZoZSULZmIR5HVf
zUvZl3GZ2RjLUPbWnjNTv4dm3R7p9GfFUgY1i4OZor5ptHIEnZp+z4Tfu4rzcv4Ocoarp3xUWIdp
VsvCizWC9wxlGQ07NavRci72h9YzPFWZrSSHiCUx4ELu5VrIW4m8TSKGO+pPdB9VTf32+u4hGhcC
BZ4xn76xnkdd4KXAF0QaPRynqHyMZBgKMSE5TPdtesGjUexaFg34UPMZWJoA43tbQu+p3VQwHrmr
RD7qT0bOBjrU86b80btnCtju6Nbpt4gE5W/3AwAeZD497+dZ8HIkkrWLZX0FrRSHv1rdq4R6VkWE
tP2xMcozleHQvS1CCwazsHDCkiIGx7nbkHCCt899WR4iD2sMVmxhe5xaCYH7JJ78BfSHlP5eMRYI
Hcx/35no5cPpkyC5dtIoA0V6DwI/uAVmMRUoChjkgcKtfzVe+qDv90H9LXgJ3k0uTdO7BDJqpJTw
/ThXCY/ldhVpcUovJ6sle57tyZnl76MzU4nvlcmNkL0ms8YtLIaSV+WPWlia5T1/7F7fyXF1DRy8
p/obNEnwEnLrgQBfVu2ZkEMyGnQ58Zgof8e2GycWcoJBHQEID/sSn6MMLRod6Du9A3B7vccOIGob
zkOZRjeS6flrAEgukxP8LUdliJhae35dQCerfehHV11XxdkZajdAhyipRTpF2QTbecw6rJzMvTMM
OYr9FInFkEcfjFGwBMOe10gorpHdjtZtlQ7ANlIjXBBmkf9Qu4fFlK2lXjecn0pcA0U+kh3eriAw
LduJVO7HGkMfiSf+T1clg4GQCJI66OviWkYVXpQtKjZGPjbgs5qYATDMy1G/FuWN158wIh4Xzrhv
enH9gi3D7uYBz2M8naDQjJ3WGSyZFToRXMeUYGGE/u/6QU2wy+NZHPwzY1lboitZ/xY3S+zT6h7V
1aAEaS3xS4gUL/jZQwq1sQXAohBgB0oX63nF9P/4IaDC/xkOflERMYqe1RvOm+yaMtnRWiCLDd99
LO63WcfWi7S3C8f3b2oNvsWm0qmXbYOc0t7uhDtDA/JxaqNb+/SFYvxfvQlDFlHv4VvK+TSPahes
Nf9C0mawkbWfIHUWG+JkIgoXyCpxrDjPRLHKvZVgZM3Q79KNhk0H3CIV+mT/5OXvhtqA+FyC4HYy
Qha/uHEFEZLdOTP8k1XtTH/BnjtFqZIv2LXBCpQy0IAxS48RadbURUUu+Na3dqu/4v8uv4tLN+WK
1hzgpchLxib0ZnN++P22TbERk5q+ZPzjO02toaNz63ymmyjtpL6MK+UGjfe37V6gr7d7Vv2RYF19
it50hA/kD9azinsQdoLO14CThw+fQaTq2o4fndapKNt2b2qN1lpALDWAEouef3bulbywaeb4jCVS
y+BVq4zZzBUYl8wimC+f2x5vv+VN/L4LvagPecDyEfKy8hTw6bWs1os7rSef1PWcZ91VTZKfhohX
ZdgLto6RZxYk67tz1fhwApOUkLO/pY0TlUbaoQ9339OvXY6rVzCW2HFQEE9fnDUUt+eEbI9nEXw5
j/sejHWBQ5bwlS4cr04mKWtMUT5xL+vp6C+ahlUgS4Pilqf1yxIIQDPr+3RUTxMT2hgP+EkhIsv2
2aMQS18UOt0toVVDfczU/MVDgddnFhd5i9tYAmhcM73zUmJp4FAyoPaLmKIoT3UQu3xLxn6m4HGg
LtGCZQKnelPUaQSVqVInqxSW2LJjO0Fgu8N+o5rf7VwB8BEoAl9JckOKdYaVEGMcErDu2oDhNv/X
9WPyV2sgn+E5NIKAiowAr1kb4tgpQZK4oSGQWzxSeKR3sdkHIpzdb5pE+q3Sa4WVdZc6YzSRCYEJ
tLFtou1kDw2na+yUK6axtAK86kaPf5pc6a5vllwEF5VcdEVInsIJO4I1Wcql5XsoW3Ey7E60Y3aO
xJqgBf5cwQOMySJQH7GwLZF7/J8Wnz7I4TmCsevFi965XeZemmunWR/D4Fx1ZrmFVYKyO9N3Bs60
q5LYiGj8TriBe1GfiHJA6vYpx7appQp4KQ38IMj9sywJGmn8uf1/nzMRzNy9Ke8nWKAIbs89lmkU
9nV+D0Pgs9IAhmPvPqgZyTDSxLg5cekc9OrVMEgfBrVEjg1SSuzog1eTJM2UK7NkUBqvIUef1TMq
uP/htmspSWaU+FW90EruPS7abCW9szZIcvGXK7q2Ms343F83HchEJ6sDCGUfefT+jnw2inKdVUwE
9YO9W1e4paiiIuXSavA5pb3+X78/I2njvVIK9k5x86AXXs5o1vHmNWl8Z/iOhmuyCkMtmY0YMHyp
4JXObZK3f7osxHfABgOpKILpICFrqJ33Fyy0IiJ0a6YPv1EnVDaDhPLO501ej/YwXFeaokbv7tCr
EYlILgIXe3wTYkPdKCax3hAb7iazuiee6MgbIhDWy23Bi/Lb3nT/ygKvPePB659gTTU0LGi/3KtJ
N7TACkO5i+xC8hA4BHXXlOMMHsdKIGXNTqw55GqAa6qJGqjXfAS6FjUwdmh+AwjorRTzkmA17+LJ
hCBD2UOJSw2uP35yufZ8OlrNMLUOWXPNJo5SdnfAthCll+2HPXqFjhyFTfhN9GrLXAG6kj+VhmEC
qnjxUoVlqiZP/1tgAozFGQBScB2TitkqlEe/zpgOjraLKOi3MYxkcGcqUN0mlefvCi3wCaLWSHWQ
5u6YzXfjCLb2ukX3FYHsO6M6Y5J6d91+k2/DVIT6PplFXWJ+tke0bL6jcfJnk0qE5VODunSylpFu
LBVXnSCrs3Fjs79QYWEC6nXxv5z6YMZVS4mLiemt/kxVR4m/mUKKjUToI8YtTPEdDi8Ek9PdLihT
LplSReJMtm3AcMfNfOg1oP8g4c+UMR0TMkhiieil498I0fW1wYFAO28+Hqg02udNOMxqMpTsn953
5WyWQDEiicTUfDWUh+ZWcuGAaxAqQ3n7rmSDSpKChiu2FNXiC57QSts52otS23pQgpONoBOLxJXz
YXUcZI0ALXXMDILWRDNZkAUWMQ8rqkJCqJLVlkQbHAvDR104jvYHuu0K0xm4/5wHzdv7IAYtfgSX
8WqmbanydR+WSLvnOsC0NZ8h9Ujw0jg0O2nJ/rP9m5qCqtzjSyv33FjOFr8Nnvxb4l90jmDHejWq
i+dkp7wm6bAOGdOf4iaKih4BLPVQjY+s7qs+FJDmdVIM5AZ2UkmNBNfnO8J6y0Ux/dhVGkC+vv2F
C1yVSm6Qva0fYf3ipH0AA//X+EDE54vrsKojsEHZ3oiuhrCf64+kx05rPWiRvF/6PnYT8VhyjbIA
zexBvGts5AkVUX82xpJN7+BZLxRoPpikJ1ANyJ6hSskWQxO063AhdCPY4n6c8ZpiTOaoaYKv8l4K
vnJzSU3Tk+DN5IKWzhMXpoVIOEQ7Qs9VIhXAH3KDeJmDT0LwlX+JxvGIZC4byDjzj0ztjgkmmcUX
LOXvEytYRWF3ZRmQftD0gOPUdMQFLhvcP0+xtZ/MYAuu8cqFJ7hmTTwaFhizqUPblE2eb32iYb+2
E5Rj0L3EWNHbCET0uhxlgBXPMl43eL19BQCCwDky+18o8muOxRhQndIqSL9z9WC81Sl4dsh9t9mc
7ypC+p5+fW46HdzYQSbYPQV/cipf4MyQLi/YuQPwpwrfjIe6QTlm0Alq0fc5Vj6pgmFum/2WVe71
3dvdQdAYycVo3o7ENOp6BUp+UeUSTHZl5tOgO2C/JmWba01LPttaOigxjkNk5G4ovOUYRSiEcRzl
gbmFJGXUFxwBg5h9haZbMv2aPk+/LMZ5b14q59DJY1z3w379TY3lzJ1PbJ9688367lT+To0B9iv5
0NPzUEjkpJxtPy8ANb/aC2d3Op4DQvWl5JiZMY5voTlTwoiRRQlmacThXSnm42j1jap6z/5CCtk6
Cg0+IC8YSGJdpwATvGiKc10m69ysgZulXm8lX0ELBtkFHRJNVApBfzMaL/7krluP86yO7bRGfOof
9FIN0dibHddYsCSbBtkuCwrEko6YS0rC74ICLCORJBrEN3xpDxwgIuT4LULdZmelzETbKfygerL7
ANk25T9i8GuyeoAZmwt+D36NM08Xr1mmoD2WsM5ygH7qTHfIxnm6ZdLoq7dqjsj0scfw0SmDCsZw
25jRaYpV8NLI+YoNzdBENoh532mOPvToXVFBFJn/TmTKYnQ5NXtYdNcy2DoCCwRYQ1e/X1yUaALE
oKX8nGdfb1449cfbvVAR0oRWZOggmFcHVuJmeF1RTAcsgu/+OQf7w1LBztpBh88CtGBE8gSubxiN
+Is/yNPfNSZWUTvUqHZjvqQTSn2Os1GydwkcmofIQt6wkqSOmqZuMK0xkY0IGQxeCIbTBY0FZyg1
8FmMN/K54urPVYgZwf6b0MG8HXEBz2g9OSx76dQ4+yRY/7qccDzRp9xWmzp+STcqKVF1InZ62wDG
veMi9SUzCscJDfgV8YAPD8+fR4RLs9sFNWGhsU902e2YdiD9SFh13YpC3wimziXmihZVa+8AqEUU
g9223wAanaW5E/rgL63Vk6oVvPje2v1wOU0bavU9tEbBez3u+peIGNy8PelDACk+GelTjRtQs00m
A8i8DjfkJt/eX+/Xo18PkDgDZzeIlqiIW6313yGCJTCXYrLi0TN1PNLjF/5jrFJjBfPmk4hAknka
1wHVENZscul9OXJFQB5q83/+ERN2EvvWxEKtWppRfE6YICHw/iUc4GJJk0koSsh2PFFzdoawXBL7
S5RS2m2AudbeIt3OXZPjR8UkVusAb/TEjKwumiaNBNcCkQH0VbpZEuFrZpl/tXfnrHjKiqOPUtpQ
VyWGrTWwnmrrQWcp4PQYpwSXcbMc3wHZGcZ9aq/R+bKND8pKjHaHdlWH6DF556rYn2BUZia8+U9i
dHjZAvpNh5bGQ+QiMBH8MO2zDll3KBJsL2eVjC0eXuYpLGNxZLMQ8aLW++4df8XEwYcOGs/+ZDNj
XRY2+LSZ7sbg6KU5ilPUlrWvPcYcTESt2GNTIckzmhD3F0YfxYLiqNT7UQz9uG+Ovyn9N3Dg/rtX
rtfFdjIF9ZpXPLeYlEoArxV6KdDJ9H488hZRJCkvnnDjIjnuxzI1dOxuWVlzj4y4HzqTkfiRdec6
NW2V1CR0CRZQ2fWhMdf5y6fuZ9Yqq4RSw+V4+MRGrNJOALKrXTRNjf8SkbqN25lBmuq54agqYnxL
ebWDuCNoipcWHy5g4b6Uf824mEiDnGXo2fv00JpaIRIGtwN3vQs3bVxcTNcQS2M1vS0ILsgrjbnB
C19FukfC16hym3TXhzXHrtVM2C9ZVoCuNwX7YhzptB7h0EN3yN1FCtWRVew6Vc0rhm/8IIrFa9jT
HHI3vr/02EXIMUecvtDo70nXlJmeBH1PFcKf08I1y5BSAPNRLGFyTn1bolccCthaDiVghJM6LHvm
NqUYSphr774Lo1nXnGy+oRyu6GaJf8ns/C3EblldGRroZq3ETfa5dG2O2dr0iNUBtQGljTDx03dp
K+7BPy3dqnicgauiMR9qYYJrkOfS07ZTOUPxER+iQ4uJ5Z2igBz0d8vbQoBoKXC74KkrqbFwTDrj
eemM1EM9WmN4geTwVikMxngaKQc3mFyGv2M6g4glojkn87AiAhu6/g7eJkIkAIpViVfeD4bzsM4v
ZrpTdckK/mSX2U3EnkSqKwl0m7yCS0jtcT6sBb1gIRs5V33jAqZs5FW6sLp9d8r3Qav7o7UBc+ra
DDIBIH4ffqDoVk06lwaymbtgFSolHukRPXNy7zNcnwn9bnX7tMcDHidsWiZaYY+RrNcTig89Sf9u
cAXQAu/g7X2XbrSksG1j1P0+AtIeG5wFQzAaps0AdtDP4SSjXUoPnHDdNFfdDR10rBTDOBSMGyho
gGregkSu8YJHx9VfnrW3+RzuLO0v3qeB96uc0Kr9MAmtMLOUq99rqzm2vo6Xf+aZTfVmGb482IwA
XCmY6xsb8I87W2qW4kLlEdfb9/esJKxDnXOsac+38ZaN9uLssUHr/TBXulZ/Lj6k2deFwV1rRCWC
Rhle2QFI5dwosPqvuDJ/yo2vmggwRaTkC9U97E6eSAdpZFBXPtYbytu52i5AUHDmRvyRFvRpxu2d
G1YwTRPMblviZfUWfbeFU/jL/lZt0/zileKnK3H+tfIgSRAmF+t1oe99Ix+o3EC987lYoKi4Q8gl
msIpJ2pGx9CAX8xVhuflXwHrrmoYI/3WjXlvW57wJmHKmua/7Rd5qoaj21qwDHz3fYMtwkdVlCx/
yJTUlRxLUS/hfnEfJJkBzC/MCKdyypbqml2ExN1W7ARvG01eNSRuWy+yTinGeNpu+TaiavO34/2H
eT2PpxSoawDZgDXrOIxGtH6sHJgaZV26fdO41AXqvKQ4PUXRKhxfJ8yqFp5Vf3cBBVwigsHn0Ov2
mhnFsdmGJ5Ie/ISmK/8Cs5SHLreSY/ctX8qHcgcUme8GPOUd75cq6HZ1j9+fN+ZE2Jn6bZcWJ6me
X9Ok3C1miKUCdE9BKyAqyprKsa9agjGH8DPv1zWWd3+P6I7VIJnNxsHcR73SeTwDXFP6pkySV80H
icKxPzNaXEruq1AfrWzMDMd2lSrAm6mm/ZPYIfxRd1t8Fz+u127DV+janazNZNHnZwwbQIMBG4tQ
z6z7QREHRmFKl2XRd8RaKOvFPlUmTPqGxpyW6gSy1MzTchOAJ+thYsexchq7Yk3OlrHLHFIy+Nhm
Y9rczy7W/LJ+iGAe7j40L4CLS7XKAtnyd1VTjV9bsil5qQrFduEprLiIYWbp8X4wzbOn0Q1oHWsR
n8JFmPdvXi9UACNcDBpLtX8n8BMTt08+Nk9XgISHVfZyXLY5rV3/ZlUC6PkvyIvVWAVjxU8V54B/
OiVBaSGlG6hLd1uME/floK2Cz5KlcVFBxFrjU3bmrWVYlZQHeMtwxlfCJWSApUxQFY/GPolRWKDW
dKCNR+NQwLddwwayyKsuf2S2nzzJ3F868jmIgiGuYoBw3/HW1kChhDSHZI2HTjWKy/dmixHT777A
noD9DggW3fvRfuh3X5v5UfDM7qmkaxpGv2Tst//MW7/y4EgtXxCAuO1gttUHfSFCNFLiP0hkppDA
X3w/RMTv/D8fuLWIbagIndF7olUZNfpoBsKeN4ykPmHKKBl6cVlI4h3nezyO7RzSWVR5SmNYiXA5
/3sXOSW+x1e5X+YH9Pg7qTXwRcWMNO6v80ZcFkhll7Y/t648EzncebnZGZyMyif/D0xxhp4bF/tE
VuthYz4qSygsi+Zs0iGhl7DlQZ68QXxCiTvrAyEfQheWK870SLSUQmA0gLHANozrqNy23Y2+bZ5H
fpYDXvKehXOHvM9bjzIlMoyDzkmW6DTNaMDuMVl0gJI9mAdYMoP8UmDKDGzbxN9euSsA4b9ZlZgA
ukovXb1waXfZW15fhYRslKYGHKmQdxOnS7Iun0X4Tcix7Bz2XhIy7RcjpE7ljMBDdVxfZiqUWyrF
CnvIx7e3kd8J14G5Va4KnM+ATrBPSK7iaUHGXDhvtuoiDNGJXfFTHiymd5X9hnpzblTvAHbc/pEq
kNIOjeMV4Gqu9gYIES/1apgv4V7RgHwAudsTlNO2api1OpxUnTRpzjGr21HSLLZKtyi+RYrPdLgh
d8tZaJyTgaqMH3V3CeyW0xWSvt6SsoHUjyYJtv00svlFddxu8AceYGZVfzK2pLmjBH5TwzBGTwqt
DSLYgANXOHOGyxro+mXhAkAzgZpsbSuDezeCCSinLNN6bVzmKzOxOLdsuEGnUGXNuxA6ZQzzU9d9
DIdk77AUJtJK40sdkXmBZe2tkvWTG8j3kOMWtQhijYjwpFz81aZYZJfWMKibaXqWt+tMSamfwXQH
XnvZ3BxiLh4HVcs963rISKTcj0JC1O+fjROVDeWXXEC1Dm8IfWlJzCWJxNLatkUqIbFEMug+GeoW
F5Z70el6UN36hMVS+VSlkozdX6WclK0AVRLVT7yaDv+mEMP1lzBlLcA6yBO0hZO/IsytriYMVdAT
yUIu9KF0I39FjBeHHLnmP1QuUhArzWZHUwNcpNIsZadHT6luHDztBEk09qz3zbjHOv2VdffN+BMg
myaq7nfsnQBjikiQ8TwxnI40SIquWlMAaz1ZI+oP8qXbaft/LivGHOTHxZM1sY97xkdlJISKRDOv
ltFQWEZJQ+QLvft9+N6dLgKHOTDUc7j4OTUk4Gxkm3nrqOlNBUAgpy2xQZuZqGDV39igDIcRZ08M
pNZ4pAGXjgl0kwsAu1j5VZHZDqj/Fg6DzEM1mhVXF/W9gazmV2MU8lErKxK7SllcGvkXnXvrAP49
3CtqJ8Od8Mt/CcTMdt1oF1QkBl1VMW2RSVO3Wq8Wr+bkNSfqnVvLiFHoicGIZ9p4FjjYAlbej4CR
zAC0PKC1Zq6Wei0g1MRBo3QR0XU1f/uPcMiEOxfYxlQ0cjx9rwa1c+kNAP+hP9Wv9DNUxTNRCsV9
5xXP3+m1DOn1KEjVoQ8nMouuX8O+tF6C1Tb1IQwPbybh4aMuZcgT9Mv+tro0KYr1kiDZeFl7fwYh
V7hh+mUguJT7sbgRfxg6820aMOIbYHrXug/vqWoo46FGJGgeB48t0vjqglHPx+U+W5n+UntQiGtG
9B9tYQ203CHbYRI6kQVzMA3Bccs/jRdSO6pbCxlBXFfBRZFsW4+aXrcISBI0c8QWsPeokLYBY7L9
+MJ3cC0giRIV6AT5zaMcuEhcc/jspmKOUWvAaqgvSuo9UDhlfVdZKIByFZoBx0w0ns1/CGcSJm21
q0BumJLedaqTYndQcnEMaNvYa0zLoC/fb4sFT0VFL3Os5Bzk/cKy4Xea9osK422Ar5376usrxYAN
dfTphxncB5bBM/TozXxOBhOHpRfEj8QsFRxhRP9k3CbfRV5/ErAmq804yFAdiBIJHbv5qxLmctML
G99SaOJRwS4BCHIL7WgS4rsVH97epaK8oLj9u+pg/82V7E62791418L8arng3sLiffJhRBcwwihX
fbPArLYD9++6+Wo2E7RJ810k/Jg5o8K4rsYbcUH1yMTUFJ8F6tHmonHHdoSYsQm1lDSxcAy+4K2K
zkwxTmmB5OUV3DuLlZRMzU4YxJKx1rfTac7bc7ZKUY0j2CJ6n2XBQRn7kkgKpVqqQxB2xHykocsS
tm3d+A5YWK9igZ3t1ovj8OysDiXACzc9gTU7zlXuLrCS2WbB6QkbjeBzKFUljqM3og944n6IMixB
ErxZkW/JA6rbOe2xca2UsfI0+tS9LEOuQrp7kywv5pE/CzvZQdYUDv2/kOqPcBBuy1wLXs7RgTTV
E+cm0O2CuK7g4RuP8sPJFGBgwieQmI4dpJ8DrbylROhxZy+fmx/OMuaUdgyWmEx3afzGMwrFbjQd
Fya9BR2hDDiGsTzhbBlYgB5+bVa/hN7QB8BAbVkLGOhUr7mnUIFRZNBw9MmHBSyzPyyFCK2qAexG
1KrpN4sfpxfP9r/USrWNuwHlum7j0gWrAUdstNSSnMTfmh+K1jpwa5SzCeV/NUs1ILeFs587F/zi
4OsWWazM1fpojeYhZUNaYji75Kikc5vmjIeOXRpwZHwNeWQp/CxMstHu2DmUxJnGHL17MRkLQGbA
Azu26sevM7dogwFqJR04Evj0Iw0u20Z1vjWIY4J/e2fEmjN/UyYbE00LxUgpOm0tunOTiID+1WsD
67nzfABkI0SYVKQNezkterxEQWufxxKnkL5JfDef0Sm+sXFSHi1lxJuvrNRKoZ4GDwDkQPKo6XOf
sqkugI7vdnGTt82lCTDQZfhqIcD32QwgDvJekT8TdT8eIQbIrunbXYrr1vWzjk/bf6VOjiR6MjcK
Xa+5FFN9Kja8XOvveJQtT/fPX+HoUf0akLGno00s7A8d2pAXsffDL/iWwJZQzU9tUQ0n0voYeUss
VBQr+PA6OPWWAvEn2/Zv009KhFEwm1A1SRaUT1ax7OrblTOq8FEboKN7MxF/SbGKoUjgf3XABvVZ
oGfnsEj0ri/2MpYTKLlwhAlQhaOTBpQBkTQrdLBAZ8c10npfaYRm5ws09imKbXHg8iJFXGltYcdO
lw6KRuXReYbM5lTvGeNaL/IwH+OU1OW+xKjPgn/nXXgz1wue92Xf6uXNohzQZxoSK7/zdk1qn1vx
0/yYh4swxqejFRONcIYnYswiL96tY1Py+TqF0SQOuso5EPexszy0/tcusdgyJjb3+LGSduf8h75o
tfiixBsVTkmM/BT5lT4oe1r6KuxBV6R6LxoVtDxu8ENYgCULJL1e3y4pGUsM0ZZv6cVnzag8VJA3
ha2p94/O5OZb6gpEJWrmEBLt5flQ/CJBILJiaRSjAWYu6+DTP3eCa7fyWR/Iqhtp3SW7T30Hma13
WCyGVLDIu311j67pFp/WaZyoKg1+ygD9nfPWItBaQ9BCtGGPe/nW8G//EAV+0r6e9eEcCpX93M3P
cnnpZY4urGMfEEDlksIw6faD+9gbUsXyVuMB8H4oCseshMLlws78F7kOwe8hE1b/uGoOuP8MY8ab
MNEa2lTDex69PRdh25tQI5KLfKkkcIJG67BcXqazOuKHsEg0NNuE7hMBONKm8Lqv4OAcRSnB3mH/
JkdMrwJ2yfUx3GAhx+Z2jGgTOmMJMGcvGSz7TKySfAEc9ju4epqyoSOHoCRLnwoSZ8Dq98E0FHka
q697OoOuC1qJEO8MDcm21sP+F95mMAbxL9CegCc/S7NbA7OhceLAvIDc1wv/L600tlZ+5XXQZxI4
lYsVVe2YdQvapvuX+OKnPGVm7tE8eK/fzyt1tHipBI8SX7/KBdEyGgGEWekDu+dBznrC8M5hmB83
uYuE+Gmyu2uZcJH8kI7xZ/ZPVUle35OKk40HgM64wTAKd0TUpm9osUOjQsNxbV6Ju4U02+a1Qj8K
c6Cwrc1pfjOb4DYZqHpDm/hm8dna5+K3bru7w4lhDoJVuYX0AMbhoY+DtCzuD39Qir27zYuUquhs
qCr4GcMkyDHwpMsYiQ2UFTFgO+95zWsyXifFAs9OB3XKp9ET/fAyqHQTqXc8SSjUxRMSGGHWagTf
9dNAfperbu6ch+VzsWmTW/i+a9EbMlJfNYO7arX5WTbVu1H6JG+tJJjn31hNXSuN5KjDL6lSPi49
PWUq0eXC9O5GnHwo9ECUspgQzyhGtirGDRDMVlwMc52swNrvoE0tpeHJhrYNY8PMBxycqcpdMkJw
C5bZoF99b5sznsTvrSDh/uZR5D+uN+ZREHSxZl095VnqjUGrc9RRQLltCHv1WJf9mhZuDGUHWMrs
+s874jLC04EF2E1qAd7sdtiTf/5jzwbr7ccGllBnYCmUdr+eXhwOCqw+ePD9/med59rAoeDGzv6N
pu3gg/geFkmIFpxsXcLDFZOx/81XRAm+DzHFjv8uLZ/D0xx0mcaDvdRFcYERQ/eerJglNsTgF7lE
hk6ZzNqmSk3k+3z7k8Vi75I0VxDnBmqDdCdKekriRi1VP4LVnXI0I0P8tng+aQxLWrVsrzM2Ks42
9dNshJLAjKydfnF5o9EtcxTy25FuDeNZH23E1mUOUSLSyCD/PlF8KouZbul+GYhkgq8ODkjRSpVz
XGpblQqSKDSPv10EIdojJNwRMusFKax/mvR1d1r60zWxUqDn5hQ4aiWb2TBC5n0yszvwTEbeCG+1
EW2o56cWlgfMrlK3OKKlnM/PYSNiPjnykFGtUh+4ew6vRdnmM9ZKfKA9vr9RDWIhAk4mqDWct5b2
mqSJDk2feHAlftVgDWbs8uypSo3vRR9ujJMc1j+E5SIRNomKNcTeoQwsQrbgdWyl2lOWhkPvEj7+
xppvXk4xFD/ixCWgTmnjoaQbm2xJi9UdJQsSI0VlINcitKfCutAN0hl82fESdI5xHxP+8vxKKTHE
mtuX0vNlkiNU4KFPAgumuC4TbpKn1AfG8C35wRNgLdkpsoHzUHWxwX5G/mH4uO4x+rFcLPSQEk8q
wvpjVf5k91p5zk80U+PGHneOWUcDNdVGSBO17W9rVxcthsVGhr72/J4+V1IF11u6HJuDqH6eNft5
/bg7rkvO3WaYvGJLfpD4nDdX3Ow9EqoyDW64GAQHAf69F8RGVSpm11edUO2SDxKQOJtPwbbKpcmj
BQ9E8hD31OPJGBdiEtTEcOzUZI1DDQ2c6emo49IG5h0xMkyY1RSuikeYqFrcPY+DCeTY3B0yrZVX
wfV02cP/ztc1GMXoegD85M1XRaIIBm2JVfGS+F1uj72CTCY5Xo1wF5WIkNG7ndDVQwDxKZha76Vr
8Gq4/76MqNhdcovp+foFnf1CvCzK7YsUdsZXDCVK3HxM6k1fqwDuqsj2RwptJL48IjXWQuuhh1hd
VFjdre1H4lfOTQF0xre3rAlYdHyTQQdL3RNpyj/BVda2m1PXcVG17gsU30t3e9iTtrSpNmXW7ArX
8g7dX4iC8H1zs+YaDZX1siSEoDh7n94LWfwDFUW1GcGUyqNOTqFeg7WmbCaq1SAck1rHZevHw2dQ
TIj4Xz88UoHuzBVUo/FWB1lgfSdgk9k8aUXGpdXETN+Njs/+pWcgrbO8jt3houJ/xXcsk4D9GD7J
rHCo3WdT0lvbLEqA7ZK8JLyoCYX1YfhSwNFUU5WGp30X5zVdx7dOLgT+YbAlA+5l0zcf9BOn/fGa
L8dWXKSq3eypU1v3/bIFEOBBRi9xN6LEsdNSLo22rFPiIg6bLoRFB49hM+Iym7uFAadBaw7ymVUn
qBlyeVXRdd6TYOFEFBv6JIWggVVFsqTNBe67vbgfk2kHvS8Mdw67c5bGOwY/qQUiDLqaq52YhDeS
6L/vEagqsCM1XctvzoTELGiOwall1Cq+vvIMxDWKzL/a42vGeBqY+XFZtYVPGpBxHuSiJIzLolRf
pFPI/QhWe6oSMzUB+RdiKf/Q12AYiRZeW6z94J6GI9kfQeez75+73c6rGb1OMIBm5DohddrlEz5z
IIZlO2IuKXWVZpAqff3nKwOUrO1bM80DLC7lhmWMCbNwXh6iUfvJRXt8Hq6jRJ+dgA8KDrKKtfPI
W0XoGExcXvsS5JJckyfBLmAhUdZddS92au1TgX7L6/51DWV0vQea0fRAey12Eh7cFsz4sxHy3+ek
3K9Rwd61Fpeh71ZrUKVpJ+TQ03xdjEC+myeGWLGrKNAf1zlPMASG7DuLiY5urJWB90EDhG4Kh5lA
7o6TI+3XkSI7LL0aWfCgWYF9jLZMG+StQosnjec/pT8AQ8ivUVXVpTL3R+nZkMtcDC6b+goUvC7l
zJ3swqjvbispKKtFttEHm3/JvMyHaqoCcwWEVb30MJOigbbw+99qsW7z7UUPHIFGriquz5UgU7eK
3Kx9eWRmNwHVJ+ktvQYN+P7edkJ+N4xDg+ELwo7V31N0FcQpAsZEkfhLLGE5Nt6jZAQosCSys3Mt
bKMSKs+dD5LV+UhDutQiIP/8RD6R3aSdmFMtke8mp/w0HP5tonfT0fgJ5xIdUr93dXZvICDU4TYy
bDzRUtm08M1ANvYOHYKIk43r3p5AVrJ1wuzGQ+zB5IbuUB4LQS5WDEw7FK4O9R3GuoRa0sRydl2q
oiUHGhVckaH/SvokfmKPOlWV69TdV3yKFY9HL70j4n+uRYD3Yl50KbVQxOPM0Mir/fFyWre4KbT+
pAVkH1unBHdixwSrNAkHjUyjqSTlp8qb6s3s3XFPl8YvISqEdTb+fMPYydGsqLzfKDyQYrGVYoec
CYhS1QCZMrTfAQ4D20+ye8dOSYAgjNCUq3WAY5niKlosCsE5ID/K+TZS6GyL8k+lrDXdTRCDu0jI
doqql5JktDzvft0nOYQbUER9G3fxAk7zb/IoT7zuOewbvHcnEkJyzBqr2TCyxs3sUJP1XArOealh
fqs6G720RU2gFTFvL0aaVH7q3tNWyDIASq/8TjK2Oh7SCBHhNnqC8yit3sejySsgksy9725vwEBB
l6JgJTfWcukZtiw5yQuIX/3Ea2pdJrVk0Aq3Vh1rJZuvDVePsC6gSv7LyMg3R7sxqmIlaPEb2D+W
QIUupXHtbqDDZ8AFdZ/Jzi9P0TvlJNCexZ76jeos3phQxPpjHhB075Z94nLc9HmQ9W/zsQLM6sPn
erii/03cp9XQgMzuh0lpsMgX/Q329ahtVVKkFGzUQBSZFqo0tK/PYHGzSI7Z91S4ff8Vr0s/OC3E
TULdbsg/M/Axzxy8RGZcCWBIgX8wuM3Lo+iFSBmoB0eqNGRoeQEHi+8YAm0xCT6aoa31wL0UpBzy
GXbYOf6NIYuPKfX9iyPQfqS75yM51eNPWbR6ZsJS/ZP1gpChMYtUoS1GtU4zYSBHNhwhs8DFEWj1
7q5rXubrN5PeYE7DC6vnjsaOWZh+GjSWAErC/RlWdDMeuTSgT9UxyoztF8DJ6GZJhk5Dngug9AzY
XMI0/XB0a/is7DUSOOAZTKDllpJ/r5MkpjRNTqTrXDjX0q+BiTDQONvBCzLKBb3nPhYT51kLgzCc
lfVFO36eGR9AXiGu6ZAgwaR6l0O0qI14VvooFA+Mr3q5mPXTS91akK2igy7k2wvkFa0WgaeZF1tL
kWlO4Gnsqqtd329dsUU4QBiEu/3+GEFKoNkNm8G4kImxMav/M28gN1EaSEGnwIYNywL+d8eJ1Fdj
YyCtKGb8+nlfnsu/JUhmIEq3HmoZ5wJCrtdJSiTfJ1TA6Hn6j2y2KtNpoCiNzwMUSrS8od896k0l
xgTVcC5odIcY01caMr8wkI5JPXz7eO8eaLvs8Xc+OA99Zv+ZdSOXSB6KS03WNCnILhVY0owN1z6b
38nAW6nyh7/jqCpOqlLNkMPuSbxwprwGKfVaCFMy0aHwavxsXnNutmtQvPGMlRg0lgNXL1pldTKx
6Q7TQrhSNmfSRaB9aI21/WqNPYNDVhOWzjxs8UlAbuxvWki20D+SNDYnaCAGa9vca4TXfezoAvIq
utW5vgxa22tJiWXW2y8hZQmH+Ufhz1ysOV4aYDB2p1IDsyIX+O68n4kgYc7APT4NAbnS89/pnrbp
tuNwY9LQp/ceFFChRW8yrCQ4SYCxtNe5f5C5zOTlm8z+Al8kuRd0re/FJlrA3kvz8ufmhj6yQdW3
yS6ULHd19QGmG2Y2xSUQEaW0MKLuctIb/yxpMvzDfYwYHG7TbFSuCUPm/ovfV+Kk+o1CXuYhmdPx
NhgcnY5M+7+DIxgW1pDzw5Ye7rgDmLoU5ZawnnN+IcDf+Ykte6iNab+LXl3xbOOlV/gDnmdCYiN2
L5M9d+g6Vbuj8hnNvsFztsy5jOyMdxNzYeDHWTMIBv8NAuFQm0tLQ6tvVm7V8lbGgrohiiyCHEry
aAbdmNbr3jsjwmWILcdcaP+70eiRKPORsNlGFZ7cv6Bc9AZeGygUvjgNMOJYIOBOFBA7b86ypNZg
pXdq675H3aY+WQzNwit8HZ5/0YUNvzb+Q/hiX2g4ZK8MjRYY34dN08aGKLdvqbRABXTOmGfUP1uW
3t+suQNix4YgP5vEdvBSYYyZ7W3xiOhXd7YVE+INwHzv7GQ4kg0x6Z9IRd/MdzieCul5Elx5ARMf
wM5KBJuXVrcaqOsyquOVqwfyl5EvrQ04ru5lz8ZYDCvc3N7U4mzvR0WOgdHWpmMLEP3YZ3o2Gp0e
l5rhJLor9mcZahA7kTC9af+yBaw5WkbH+5hahkin8+kdiYKlOkJydMTgwuV1vxKypB4xNRQBavDD
on2aWaSrZzkaEkOvtVnX12pa/BN51A51TXOedv1QyMiqk7mlUYJaZ2EVoCXl5jBZZViz5R1gumjL
eYLmzzsG4a+E7Td9vscczDfGaJhWxyPhHLneCjJd1J0/NSbQ3gm/iKDnQv5bMjfNJuG9DgB5UEQT
ngG+FUzCRe9ixUzAV1bbYkXIk4MW/V6ZwSPigpOeEL+VDcLPQjfCawwTx9ra2oRnb+97ODUhC4dG
ClzybYzNdEf08EKXW4Hi7p1aDfFoX4egt/Dy51VZ+wLzvbtjNuhxgB/k9KOTUluzepyX7JMIBaBO
TA/obIPn0V6yq02dAomT0K3MiisX48TK7TGiY1VR9A2qt98U0QT6m6Q7VPq94in4BMfjFEScb2yR
qmNowC50Qbs8UF1fEo9SH918tF+Bw5VB6kAgDeoqmF1CdtoiuJgi4NTTFXwX7h94nl3eHAYR9ymK
51r9ecJgPH1roCujzgIIwEOOFd9RTxTzzGvg2qqygA7BeUNYgB9lnN7EYjieLlGxrPZ12BPcZknE
abxcu5q90HOHGoouMtzwNPbfZ14j2P2vsmKZ4WdbRYA4Jp1FJB8oI+PedLj0zwS35lg7KZMhUea9
hp9IkPAiPSgjcsrAmCeT1z1mOJ7B4dBdzAkAB7QDawloQwaZSTZvitQPq4AAjIGFvgZuax2F3LQh
CFQt5mA/HxYdLRNLTA4QXRTjehOovAx6LPIh5OhQkHKpSrSD/sQkHB4wiu/TWxhgATKqVgE/AIGE
zYRynyOKo1k1Da3WHN+Mq+5AlJM1fnKeJfYFyEfc6eNV8izbNuE1HPAMKXAvG6bs6kX77fpsM0GU
Yg6Wan3InZR+hLnPCmH1sb8LW0HfxDhLIqTBpuWnELaqXd5eIp/6fB2rrOSDkcnUjpkjkXgbbisJ
/pzVIE3KndKhHkerNxtT4JzWB62l/7r5L5DJZSAaRNY0zKmEpD2RmN3kS/Pxc62qYlIQLUIS1dmX
gA3ZVlvrMvaxkN4DEbS9UwVHEXTtIxnOo/IHUXJzSAlMslW497eg43Ka0ZoJi6xF10Hz4rdOxF84
8nN/7xRjQjfTD5ygP5p7jqIhbASsdX1QgaxgGMX2dYA6WP+/d6SlppqDjrQe8429ZuWQD+YUAl5W
oLiHL7PrMNaA8Rk9zjAGDL4WVr2VFghskFPGulY7UWaAkUqZYYb7L0Sf9bFFaR1pwaLEOb2dsF04
7lLCeCbfaNy+pGIDv1CXej7jvPv49HQpesrT7mFuiUCqE6TV7+bQPG3U02r0E/40PR5WgsOEBj6z
S3bRHMennb45397BD0iB/1cYy1P36xZI7h6tlrvvDwm2oBeVjYCHOytgQJTtKkvJqXYy2CWIQgzG
y/XlnBpan52JMcdHB3Gsc7SZoQV+K3/UbazMAQOLkSq6bKY0ns5DDB2+2BzvJAL/qDoaXm8QYlJj
fxVtHP73jsfLya+REyVt3oMepvTzNhcTl21QhXuOsD5+MtMnyCIMvwLGfRmf5kCyZfqRxgOaG7Kk
WP87FwKssKr+VSLI+dXma7A5nmjUjz22DvJBuyfIVJnyUFE3Bm0OUHE9rWGfII5fxnwfPUo3lB7X
R+2H4QMKXGyKSmbjtpnVC428gOcnLJ4s2/WUTvy9McnAH/Nj1JmxTwzCzeJA2UOrT+/uCxM2jVlP
q4l5C2Oicyo5I35kLI9RqQJGmVPQvxwyE1cqwusKHsb9au+EZHGRd/tqf0QIbG/bWPZR3hbYQoWh
H7xcTnUusQu2vjHmnlqfSWM1U4ZxHTiDCnax0JT54guImqVUGlgq/Krt7/B5jKWVuRbecdJpTtTQ
aCXQlU8oDj6AU2l8sFWBY718J/zoDiHN40f0ms2G+FE8dCsUE+afL96DDnQm6NJvd599fNHZph3x
CjUxeOaBVIbRTGqap+lh0sPccv5nJmhPcfBaUnlY/eZC2yacQ2fysBBXBFMLG5Ebi3kzIlIB6nUp
XVOrJeuQ6TwVhxfPiy5cLThfLqSocPvt2Fu5Hbmqc3uYNFQa+hSUfYtp4xBVVue2mW44+zzWrRRM
ieAHlfvap4N4Qz84xBQ3famqYGpkBy4JzdNTERedCist44RewAbiUXORNJzxBi382x6iGjcYJQP2
56f1GqoxmY9AtxtcFUhB93pVNQUuEtkCfbuFG3Qj8jm9rpJFAS1B2wcRMfsI92q6/OcRfrvkr0qm
vAmijzuWuw16zRp+wIYxILDDY80eA8TQLQn4ULEwPGx64ywlS/HzPEsnYoDmV36a0ilVG6A0l5MN
Juij3DWBRlqQdaRo4CSKwChriQtnZeWL/LP7/UOsPR2ZR76zqGXNMWmp4y+1nY09ncX3vkyQjO70
04ecWoyL51VR9epqVIMqIPst5vZvjqMA5Flbxf1AQ8sGmqKS4Xxpyv4lwkgTbWIbb5Og/ADTkmlY
GW1VaMHyLc9EyrlFXksG5v0XGA3fwvmR5Pst11Dr9S9N6fvr7s83c7GI2KwL9FjjvS3Y1dtJHZYU
HZ+ZHkf8h+eoznMuVQ3wf9aEnhxzHSHe3tgQ6S0xrtLs545leFANFgb/zVHwjdCNQkkE79lw6WhG
GesLF/5qq5ZeGEfEzA/pSZikF02B1m67VXaJoJ7YkbYuQ7Br4f+GfmnpgL+S/FHHQfs2RraCGxuP
xZp/G/rchHs95GuqEfWhv0N/Lxvkngh1xAaWqSfOKYZZtvZ51I3Fm88LQl8CSDOkIFGRBCb30Ik+
x/FkhX8bm+v2tPgSMt2lSu1061vxEvOIhl6T8bTQGQPPXoz0c0IyF8wCaPZSQl5KPxPKRsoPQd3e
1OaDW00XHLjEmLJwD8KprsQBEv0XqC9IwtHUoxfHxH8qHl8V2mPQ/+6MB4vTHCiyblG3fIfFyJRW
CtXVBdjloeZSDKoN5C7emU/l7sql897X/QKAUCGpZfXv99deLyUjVzLJkrxsB9iHlNbVZ12XdFQQ
Jj7DPwzwjBach8h34oFMfvF59IUpmWH1ah/bX3p2tw+LsOMVKXqlcoUGHlcIuH6nnMyfu8N2tkxQ
M3H+WJN84edReyUnc7yTRUpuJbOC4LBc7lMVVbkUTjnAGjncrS3cKryVxz1R297nYQIvxIEm1UVW
MAFjd/abbBcHGn9GupVV5xp0UM3DYHVb32ktsIhlNTYZKzPf1CkhzpkV2cz2qyc99nyxBQiBe4j8
OOTf99Gy7Q3QnL91wIGJzMf/42BkVD1JCrlM1T5afrtYyRPhu6cNIZTmKb+51vFJZe0iwOzn9JQk
4cF1hk9JDBMGPNXHlShnpOwPbNRVQKp/V6jyV+eHq0DfxgA+AmXRtUeW6g0h6ppAbQvrQCyl+euZ
K6Vsi1qHsWgFYhdYh49v+0RCh9qYooxBv7/+RozE5KGgPf41ccOsdxmbF2nxpYDjs0ajGhci7XnG
G5amipwEP2QcWwrcQj+aBWa3GJxyoujnwCQ6tgukvb5ncP4F7KYq0ooAXHdbfvWrKfCB62Idh0Yu
dFdgz05Ia9CHb2n7MpCuIy4iacO1RANwknQyzWuPpascMPCogGwGyb4APY4FgDf5x6PMKJBxpxZH
QTDyBGulShGOAVH6oLUTOKW6rOtUCrMY7srj3iWXT0BGoZ7313kDqaN+Yq+2FjC/GQxkez0CSJ+D
gg7pyey4uhn9K7nr4hXakxy5vbfhm2l2xSFURJodbo3a+fGwIVIU+5/UF3wYOUL9cScMItPjTiJL
xipHDpyVvmpiQmqvzQGcYb6oAyb2qErQ1aAUe1Zfbd0UM2dheaMdk/l8iGCiUhMcMfqygQeXFnIR
c9HitBDJUSr+8g7cq3G11msAUXIb9qcs8preBXtYDljbNYj75DJStJB0lSeiLd+n3B8pm7hyaAno
A05iFyW5rnK8SvCZePyrUoTIj5cQE61B6zSdjSFeRY4i5R473uGRIjOOW2O0W/+QJoRRwurSMsb0
3RN+3ohM5/V7/6xtJjjU+aRWyRACe+XAsONpGzGv5ArxChIXPhs6WFXjAssCprH1Q5LmbGHTdd7t
yWreSkBAOpYjZVAik4aNoBGzRMp/JKL/BM0fgiS5KZ+pD9x2jrdpO/BHNNImXmBnylbadvapW9q7
+jauA6HAUwrI23dezPIHBCe32KEnY0+x7UhRUzJKfGjQuMV+zgO02q6Oo7UQfxYvDvdkIph4mMv1
Z38DZacOgTTeBQKU7zZVcRNacxMqype+3YDphiIodXS+t9nMvvN6J3vDju6Sbgen
`protect end_protected
