-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
MtEPaX6rJj1QmgXEllW0g60HWSfz0hBj/CK8OST9hyi9MSDxD7iM9q2ZwwcMtE5cR1wmNRHnwG0b
d5SN2hxBPs2ZCBMNZR55GLewlk0llbM/hmY058zv/PHbDDlWA3KjX+7P8sw5G8NBzZs3zjBGqvSQ
i5M63PVaczwXKjtAwA0Ag36aVcVHvpt0+pl8chEGoPN0cBiY4HrMOezkOyIfqdUM0SuNlZD0iPNx
fAbbo7g8Mu6yrKmIVJbAT1E7WqnPb36X0XjACfEwv1+oRGcF/klVzxWkO6r+s7P+v0scWnP1iGf+
L1RAvEiUZ4vBdGSla5qz9Jyx+lbDDY4LJ/5uBQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3616)
`protect data_block
ZAO+36WNanGckHH8y7p+mC55w0iqJR9QrEUJAsCJ7b9e3oWnS4ChSPX/gEpHoTgGW07rEvbyT/lX
FsEP5tWdH9yhtzX9xFZX/isMwT9M3PkGq8plNnefsDtN3mzqQ9GCr0umMwAMS/amntbFobBRLK7G
Jhb4pogSbZ8YH/T1HInPk+/jZFO+8v9q2vtXEThxnq53gu5nZqg5KBj9O7J8lSSv5413NOyz/46f
fMHLy8vp0HuL+7q6y/bbxUSrieQAwirQgpYDBgRrdJnJG6IZnqjb9vdz9wi1VuwuArMrmFk1pwJS
VwNBTcwp3GBPwnwjzHWJNeARdhfOzrQGAaS5XVzyc0R4hc1SFyyYdMM/B/H+vW8ecsvZ2HKRtUdp
uo1V49FMDDqbiowhtaI8+M/wBruzKLHvMSRmnZ28ZumglEdsyi3b+kQtbxAV7Qxf8PV7xysB4qb1
2A/Ebt45pU4p+4TaJ2tfLq/6ml1TSR+c4xdqrWHON2lGSzqF/IHryCaS8oq3YGRrkPTc9J+90xjW
ILwa1wrDFNEWSV/Q1MSyNCGFo2qFLAamKeI/OKWM07EYQqhFA7c6++tRH2TXW+Jm0yEgmqiXsKii
W8lDhOJ0+7XWg6m4/ZzCK5m5zh6hbyE7TezlhtsPSmv9TUKEozZ/TgF4nwL4Va5xGUrRAvVeOj/F
nDuvam+J0dnGPPOpv3Y+EbzFV0R7mILLoGLV+1yMYsEvBSLLN0jNx0yvcaxfUyPtG99uerxOgQiE
L3/4GvC5PAeVlFw3fyN6qczJZRKvfXw5xBu7bP56QcUUpABiCmAaS8HVjjzF0uLprTLi430bBSZx
QACNMo3ThMouq+Q2KXBZxqY8t6ytvn52v0rJQpsyczSRQgmcFrR/Kcg1IZTaZA0TuHTP7ZiJbSqt
L8Sn6C1wnsrGYJQ8ui5/VsoAqMqy8Xmn7Ows/kXt4ujsDwlveYJuqES1/JNBvoVT8h+eMqEVWfua
HomtsaQcAr3d/fFI58i1VJX6Wyjuh5ap/1/GF8GzTssDwPp6kn0Rf6fuxtaCRrRt9MqtzuBZuG3d
TpywqCv2PUmDVikduvcU3yB8QPruZ7HSx64YLKT/h+JkSwJL1QtB7JuTWFXdc4U2mCHzgQoPWR5J
MIpibYtcYZ78Zx+KmE6VaAU1/s8c6yLAmoPBVHfoUPUHzEEX4OhEkAOXp/5nke0mIIlLccPNrXOi
L3jgMLjxHlcCDw/SWdNpWzJmYw99crazt67m+H+AbnzUybc41R75C7kF125/hNsAY1J7cKHSs8tO
o8q9ttB7/x7JayVubE2/O0HQeqlAgdFYfkpACpj4jtEaC50VZwMim6sObLm9JlJJTiXvNd2RXcvp
wuYIaQVN30LSocumBdHd/YkPWTKWcFhtB5NIVEJIgKiVMJ87aF/+ZKz5vcxDNEOYpOy0KMbQb6El
/Qwj+fksiWSWDzUbceoyDm0CwitL7a/OJrpZ0Mdd4J9TDCCjAr8sXxB5q99lUaKz+QJArW6CYhKQ
nsUvqxYl28LUGsyHJQAHB+as8w5ZOWhTh6qR46f5bzLCkaurYbSFiJQxXmtu3TiNq9k9WU1oGm96
jzghwRKmXZdtBeTO/dQrX2hD9Q0ccPIJb3s8AbcsY5PLZGxfPTxcUfhTcGJZADK5fBFFlPFoaWFX
4nQHF2LMrBOek6dxa9UB9tgwxvikjFb19iu5Ya1xocD6k1Tb3efWbXVaWtL6Jk8mWqwwGDtJVIS/
lKq82WF32T8xLcjj8HFdXFeL5IvQ6Jp1pmiccpJFG3wr2cnr9Hvy9cGD1YREQ45Pb5ntqS6fuWJB
tEf78+INVEOjTY0fiHtWlbCWYbtM+FkGtVgcVBO2MZ4nKP4MOM+HXKD6HML7WJ8Ap1vptPwL/6LW
jD7nGaJJjEp+MmI5zDihqKmZrFVdDr0yUZPL/dvTJsJOGjyRBHF2pgQ4HdPOExOe+PtPgriFUXF0
AGSBS7YEw3MT1fXc0pyAZjqff9APOnN0GQJp/E9gieT+AN/q4goYq5DnOz3hWC7oZPxvcmzULro/
AItB8IGs0DUf5PB3ebP1NyjgsFh+pGK6MDXYnEz7u9OCESj7kK6fNWaYkmX/Iz1Jae/xf3ttqu8Z
KFXUORHXPvHhtjYQZx2Ml2jIhbILsvbCLPR0PriNUoO7c2U5MiIyHtTSpM78wqkv1geN7f1a/i6W
4Up7+dC6Ni32l2ibuTJOg44kp1oBT4ELOig/L/Lwdfc9GlwSEINw3P1URsQh9Yg1+xsMlcVAL85U
K3MXenzuAJIOH9P+LogNbw1zyv6urkUH0qfboSrCwf4ywpMCuae5ypbrGpW1euLCmx6r94zTJfZR
TflEGaRAhM7TNiGFlgh2H3JS1i2C14ehIG+yYAop/t2+I6LGuzvMpbRIG69w2INntsFT3fezy3dS
pf5RYmvAYol4KHLLYXZ4VA3rsAoj4t3GqSYW3U0R8dIMlKUKV7ijt57JWckn0PwxNUK6GV+OgF8W
sgtsn0a+N1HPOyQYs9Htryf1X/SvkSmnGkhBuErDyTnfu5JRoUX9yqsesAfurZEVMkeUJYv0ugCp
wjm/3qo7yy7ivQ8PakN7jW10YiL/P5kZu8ai4lsbgqtbISOZCQG4SJllHcYsQCSSxRuY/Rh6KUOz
xWQKOtC5z4pGU5hOD3Yl1nbKMKO20r2TfBI2w3WcJeR3ghdCX8q7Ua+959nEp98oujIaRq2CIfhQ
JEMC3AfTeTfo8UiWlzX/aUe/tVh1gCII0dbR4LrKMkpv0IVxjXe+ik0bcT3TFzZ5wHrVom+uyE7q
91yvexk+GIl9mU1c14aQYEl6nhFVUjX6y35nLGE78CTlTb84wGnaTjZ0s6xDTnZfkvjO6j1Y9qgS
UpwNfXjAKZDwNXDBIr1EW66QXL3dsg1Hrxn2v+Fffow+mFJ0et4vk/PhChwUkR5SXTyZkAh9q4+g
AOoABP/UriCMXQtnOxwVNUrN7Sus9ztxz1cCGFmvBuBKefMCv67a7Wd3zhySMCkWarkeDAK0prOO
98UthadDQuH5kDUUIrJWcZbp35LK/GDy2C+ec2PtQxelRHBeIbgfgurTYEFoY6DHbxPyZEesw2jG
YtvF93jX+OMiabQRcLGbHeS6US5XDVscZ5oOv6oau9KZMwYt4dwvzhjYewvfArpHrUYFKBwW54lk
cLvQ9tAUcx4UkVxVqI13Cui99kkhMn9UXRpt3kUkLSrTMUsK6KKZuefeeMENsi8381Ynb9tXzGOm
M/9hFbNA5rc+KG03FrQZi1LW+liBYNBMnWEfrrf6g/1H9HsRdKVpPqW5EgmePG/3f0D+sauTAKKv
o/os/b80D2F4C4pYv8bDTlhiLzd4Byohkzc+Cf+kjVt3XblOBAFgu7E2mrryvCFtIcF0MxQd7ui4
5+ztPc/t66j2oNOeu3PRnMXdFhkTkhSEPlp8JspKaMzbe5l7qpXclzqbOJJvCYijhFXUq/i/T9PO
jIpNB2C8YuwfBMhTwpj0XOVCv20iPbRUmd9QM6ST2lEBFWR1BZQO56oQGhDLLHLZkllY8THwJbuN
nnvbEH+GDcB2JHeJ1DA2l/LCjMASbsxdost7S0Z4U+tZTn2kxF/MCOT0XjAXLzbNmvZnSmNgyTGO
leGN1IidAtcRqOy+6vP4qvgRTjieaJKdLbvjIqa+C/f5rQEEBHSDG2K+fvt+7DfdjuDf9FlX9wQE
9LPrDcUZw9yUrbMqGXjsZ7dx7WxohMEHczat6WWH+Zj5wvMBGcp0tMggx8oqN/kTd9sBNqlTabMq
70C3UOA+k4LuBEUUQZo+fUvldCdKIaBIwq8G+UIlkL/MeZg5UE1m/kAhEyKRTg9zWqgX4q5deFoX
LNFe3qCokdvXB5K/IOGjLRKx1iv9tbGCE+L47rlILgbVvnVYrd17xZonuW815sMIJpmoGpGT/B1l
79b5rO4w9FntrArXLsXgfG7Ctw1ihewGIlpWbjpO2dU27zwUKSwIy5il+2tMtJBlxYssq3y77ytt
UGos2Z21gWhXOc/lyn2Byf0Z9b9j072hsnORdioaN9Deaa1DkX31FdAVmWQta0lqTRVzLuRFfdSs
QrPEjw0WBzSxkjtbtx6KMiHxbHFe80sDyUgCqeXE5zft+uWCqA/S/fKJwW5M/HZMyshDjveEh81P
xF5hofE9Cx9l4g2WGfpfTZdb5zEWSlvPxaKla1FL+k44dO5L5Ve/0d1l2LBthABu6X+PNhfH6MiP
D5LVAtaslw5jbxoVNGKJ5RnhrnYHr4+E2cn0mgHB7ora7UKPn4fQwQrrgynCHSAVa5ugmF4q+l7Q
rJBToXd8BnlRf2L0PLtbDQtPJHZcEGt9vKHGrxqbrF/xi09ql7WE4ASopZr3W73pbmLNn0z2a/10
MP6/++43AN23V88dvLNlCk3EFrR8K6Oprk1yVnpPKPmc6omiXVwvxw/ab0bp9CbWh/qDS7S2Wp7h
IuZl1d4GyrbF65odatU43saQo6qt7YsGvvNKBEFuhVuAJ/BmW7eRhxQQCGHzmK+amt00asGcnwo5
gt8ka7gHIkEGo6ML7mhmjRojbHtNa4bsMtKKCWrZApggjkeHMwypnOAARojIRJorOzW8SKymkCTs
hNjgNYKDnSVx0CWZfK4ngOFoyU4jypistNMCNMVQSFj0NRiuXty8b7wbmjWEvG/XyYarf17BZJuP
hjnYAH96djjdwRS5j7E0j3bwnccOMp6XrehKTBelZsjsPju+xjR7b66H1/KeFVDVs04pc7QkTYaF
wS6RlD01u/NP1f2INaIetUOKK4WZKVUQrA==
`protect end_protected
