-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NVWFr0Ca0Ufbp4LPWF3voQIopWzrsNdchsg/vXelK9HL/yMrO2McxlPdr7FjzyeFRsD3g/cuS/ZJ
QJTM99Yf+inFudRtlDxEmjBhUyT5KycKmSYbyUwW1ooxiSq+D0rAjssZiFDdGSiDKW4eMdWtFKpj
PdWV+GJ3uRo2clzH2DPgB5AnR+MSu6MXGFxnlv5U+BdPI6WX8syrAeGZNdXgEK+2zF5ScpFJ1u6i
Z8HcpzcH8rqL8a1vtN6OEZLLdw1bHhE2dm65k6HtbTqnmQAlv+bmZf9goS6SpGjZqHWzl1Rmqzv2
Ronidx4jjuRhq9wpzMO0J5m7bzO7IFMplYsV/Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12384)
`protect data_block
zENwKEpQn6vx0kSVMm+KSJ/ANorJqPTEQhVp0uyRTAQdd43mUDmu0yWPBfUAfLdwbjuFBJ2xTCRv
exSyA2uTBAmfePcCrgS/1OVcf3klurHK2g71d1ivjK5cH4H/9VdGF6kTcIF3FnCaULXrQHcJqHMU
39a58B4/OrsC/JS8mWgdGPkNRFOBNlEu9jJONaX6+VyJroQ4QqBXqII/Xs1JHL+leyGHtshvuxXK
iXvFlHmJbX6jsd6LRWOt0UuWhj4oEyCHxRTvvcEhpluo9WAOm1CGpghoPLY8BadYC13eSIWNec4c
QVUW+e+7N7bCA+XyzZ4pRO0nulsjhK6CelNamQk9xxQQB+MCUPecwAyHPNf71Aiooibb18LX2tDk
2M+gxCf+g5I5oNUZvRve8Pl50+qvmRA1lVOKHZQrPdM/bMPNhdTqY4zlrXTrqmbMjNgLwmk54xtU
Mf2IGlMwfPp9BnSU7OJJBYJxxFwp0MC5GdWNqayOtpWMIXhY+jY5dvgQrsl25OsNlx3B+xW9SS1V
4cp5N7ITdJzeB/fkLZzmJuUiDkWQf4YmiCH+pm4HUiiCXHHbpw6/rhcm0LM9e/67WMuIJ5wWdDeo
dO2JqyMKODtUrHIt6tIuODNN17/aKX+a+EAnKdJWJVk8+HxgE3e8pGih7/wlKi2+aFkOV60aTM6s
LiowvQ8tp2RFaZvIbEtxqoZ6qC3bk4ZQsfQctSo14jpd/a2MoM8ctb5ZRAu5A1umgryipdI59M2l
+ePljQtt3meERzGSHFXHmtKchG59xWi3XIW7z/O3lcRthj3ycrShCHJ4cDmJzjKOyHMeG9C78oZN
wPlJUBQ89wwy+z8lxwrOgdSFjcgnXP2SledjuXXjLKKbf2WIGZuv8qzbdwHRVwaZg2j0QJ28bXCo
kZvdm6fOvUeC7PMC//fxnv/HfLAGd8qKNmFrveUgsGU6r7TvVU+ReX1DwiCJJ/LamHhidhwYiACW
xLR/pSg9pGh9z3mNzUCbhhGRgbXrFfzmI81VuDYEQXbekf9rY/+C+VJy8DEbffTE1zRdsLKL92Aj
PKbe2ujX3l9yd646FWRE3Ugmue9gI+/Ssq/dOwBWUk6pHqTbRc9jQjDcaW/ZZrEJXPmby92K2Ej1
5R5ZFJermRfSQ9w2jxoK37NVwlkZUOg0jOZPiC8HPN6rQhDsd0WQ4QUTbKT9exA7VdAPuSj0t9UG
1k0WK3G2D/rKoz4VzSb0XDki9SxDg4s5CoJfVmiICy4o4qvVTTqc/IgktSMd5Tg6Ejch1hoD2O7x
6xWHuqeOgYT7nwjAZqvMAVnSO2MQE6udMWsW25tCorYQeOORV9eRMgmdCSaCX5Jz1nAkeR1v7uGf
NYRzWVm9PwekfNNQ1jMgLh0nGr0fEbHhCb/MXpIzE5nHBzWYcSQdyjTBCRdnasyKVL/AYid2ArV8
5Ue1B3sMrbw+3wkIj45MEttoDcAsNzRHD54l19sL+8NSDWWv9I3B+Bf+Atz4SIQJVdApVyGcGZac
qERQ318kxJEyceuFs7DUHHZ3sXvlf6f7qaZ/o8TT6e8eABtlbBueTED1TuNEyJIoyzcHhFmBO8D5
Wf5gVs0y4N5gS+6yUXfMrkuiQdp3frTabsfa9MrBXgfwBOCnt8ytVKkN3fhe+71OzAOQw4VhNWtF
8+8UYp3RujPEnDMRi9JLBVraOBCDCn7O2fx7LRUtmj2DH95uXjTZjTXwBBCLXchDpMtpbu3HKvpf
hr+n1kXp2nUYoceWu1qbkKUm0goKvOFulFG/QoR27C0VP9GWxPicVfdkmogNBy1j2Z8Ud6ZHTuck
eJUUDXmxWEtVI9bLZhQydvunS3QgTgx9Vv8m6q/JQNOhNC0VSNrO3+IDetVK3w8RI0d4pWlSJcbC
GkkStQ2bm9pnxF+PCl5tHx/eZarnz/yuN2n6oSDqw0MwhdOgW9EIV6L2tbwiKTIvj7tTS9tXTZml
PG362nWsOyMjqib5NYhprwVC3hxvfNbIDTX/wAx+woPfqmt87YX7vJ66JymQD8i2dxAsWwrwzBDz
8F5cDxQpysnZl95kksWflI0mT/DGXqyEgYdwUr0tu6pZVo3NOvBQhADZ3Q++l2XZqERJyJ4xIX+4
Ho1pNIExzvvXCylAae7txJy0MGPddy2ZcqmfExd5ogFaxk8PaMJiaGYjk0Jn+TjhYXy0P0advtbP
s2us0atAwequvl+3EUAVyWjHiAG66TNvubunRZ+qQNGpxPeO5kaLZiL4cdpk4+ZHRmnIbBT1rQBa
FqHbXuIfelwUq09QCvQH9JUEHGNAdYvXzZQTEpHVlaZsOIv2cLfaG9PIydSUEyP/4D3Do1tIy0Ir
71ejBMR4uGDZfGxkOalqYan72Pgxf1VQQtn9Q+WaRW6gN6oh5as4SXTpBuqB3hW4auHaBcmNdI02
2VTTd0We2VrLkzy70hac15aYGaSyr9aUQY9ZK1b2Sq5Np/0Opk5cSjCvRO6l8+O5pkkfA3e6ZJTB
ZiXXvDUZAbdL58YVTCCIPn4LqWZxLfa5fr4v0E1ed1MhI8lE9YCP4HemS0nxXw7P4Tb/OtwojFcd
iaD9X/4hLM6ytQjhcFqxfaF/oAwxXU3dLhbI/3oXyErr0iaUOjy2daowIUn7yajADXrR66Tw+frn
VsnEJLOWxp2VaAMKFSZ45mdYs6PAUe4lf/fcf7sXB78E6I6dn+jhsbLq68QN9g9y130QxQIhkZCh
u3LnL4f4Izb6MZZc4KeFXcCf41JODK483zBrri4TCMvVfGIAFRtxEHiTOAR/WyW8fRCkuixULFRe
IUpPsnxWMLDISMLX6riSpHAmAUWtQrV2tMS+McoSkPlP8fh8OO8GRJBoICHxVSLmtTB4qfcytJac
V7t6mEbwxlHltVgb5aCkoGD+l7wIZO0Gd/c06uxPG5SiZoqbm47t9mT6XSQOOO0/IMq+jRHnml1p
IsfE3JlMsb6qwgCyKhTt/AZT5XW+bO6WDjoSqyUIGIPeu1xiPlscXpyOCzHVeUKiLm5CoqfLE2N4
CGeK46rk9y9DW6+uQk3v3zYWcUTV2xSjxCFkcZQlYV/f32yb7WRiwi1KGVxJ185BRrl8V9v/RZHQ
7RurTh8NnbRBSXybCXXcf7FCaD/0AwO+sGEpgUV1/Hhs746uOkkHnlwizPw5KlDLkonUsgYEIiRk
wObtOgjC4JOIl/2upDQGulNDkRBA/IQ5EDZBrKND57jig+fxgs64r5SyG6hBpZ30ELmvyfRqdjWo
gMWRPtflkcholwBR6eo3NRW5b1bmNEiJij6I32vUoaVyetHZ0pkdp+5s1NeekCYx0MoQQYy55uWH
HCFW8dG07eO7y+QkOil01q6NMmti0G0QkW85kHWHrdupiIudCNi2AegIrswPiS+qyd5RLZr9dSad
LX6B0YVOqB2LCL70RxS63A7K3ZcI+tP1F5URTSMbHxvmP/ReTmd/vg5kVxdPwAIpNIOpo+X9KYFF
FsJiGRuQO5h6USw+vnPTnZx8lOEZHb+d+fkCON2EcljwO4dp3PFmEKzT4BcH3uGK7rp2X7s/IvCc
J/pqkb1yAPifVbNp18OkQVOQkOIn+8PrbjWctmxKdYUBnNwsDrM5J6M4CR00u0wDSobBodKSgtuN
qvFmDQa3PMPM7WDGnxHIOaG8m6kKBF5bvvS5+RAl6kSknS3xnr7EOqr7E4s+Fwmytx7Ha19X2GS9
Pj+BHGUAvsny4s9jZr9/NkNpJLpmKPy+5dREbcC6C0WF2AQOysB+HUwcjVSEA7k5OLc8F3m0JZ/n
xwKFdgAOD2DgtlEgBtaZ7b4qLibmIVbq6uYJmBgtcW7WJPomvZjthGf4lISRBET3FO1p+eyhnn79
vQhxI9jBlCdRz5UPPePeBrs/Q8q0f4iMx4rlzBUG16IwTpVHA81CMr6ZTFU2XGe2WYaRRI6crJ8T
aUPGlyWFXfDwsnn6Jf/g8P2i8qvUjcTYIne7xAvydwvCFS9ft6UdybID8xxR/Eo+/2HvwPM2dXEc
NvKbwWyOnD0TeHzFAQbX0HQdmy1XLH7bbViGKW2Wp582oHG9aop1PAm/aOXhyCb/RUH5+7KtpzPp
wF+7sUBBiHxtpf2et5fHzlTuCaHCSIduFiQ1AVoUo9ikqWOe9e06aEi6uyOBzXU669vJSfdALZG9
/1YZx67PRm8IzwXoUgSQWrePgCvwcmffZTp5wzThcimC/1FCuV0dm63ltL19jSq4L2bUIPyIKU5a
P73eyEVGhs5tuxhNd0mO+Au5z30vzjL5Mipw0BC7MeRvWsfZtGJ9vET3L01LMrRegA24Xe2B0SMb
n0s7NBO0vBPanYamoPpDnWET25qVt8LMdFn5mjUjYg6PkxJldlhbwhy9T0SGn/W5UIEGubCnhxxw
B3et6trfzy+dnJJ6rcNX55c3qJTcYTgFrRJZNnY+8dwZ8XP7n80MWZs4ull4jcQaIOtLDSZ+vtlL
ZDBwQ9zqlWCn6McWCC5IN8GdM8nbAdreClF2aM7Wds+IanTyEpII8U6RfWoXfdHkc2Ii+koH60AT
p8OnBriehMzk4/644asXXbm66TvlZGmEgFTAqOT3qlQPB++n8MpSFjlz35L9CFtLrxx1PsD/GqbV
akfmtrqpztI2NTE9ZsAzxAkrv71AfiUhLRyJY4NcB3uIxJcPwsoV+0klsaQ/Vh+Q7Xg9TWju+Z6k
9TryDLi57k20DzAOvgvRQFTYckKV+Ecy3GwiLNRyg0FI7rAB7N5FLT6sEpRuhGukpiISLJRaI/M0
jyAy8ZqDo7OYnUFgUMxr+hdLMJWlYiLqWBoEpnRKwpQ1c2wGNg/L68ZxqTwJ66w/iRnSQ1uSnkBy
Ho71ZgGGP1Sf+NJeD64Zm9okBhMdxfbuap7Hva/8mRf5mTf0RqtzcFmM8V15vt+tL7mGSEfxx6aj
5/H3uhO01Bc33GcbQo1ueUdjumRONqGIELLNIQqfQn6awO4B0BLKC7H1NXA/OrdRAWQDohcZ8BWW
lZ66S+6ZFVtevWfmHdFU6LwpH2Se7+IYIjNG0vNxoDEdYegw9sx9gsMMXJQnZMwRlUk7KR4h9Fna
6fKteSLEEA0ahn6qLFWCbGKN+7DJbiiFdhtXh1eb7i+JuR0u3yrscARqdOSDL+nYPmpfaP3UllYP
vlgTRetEEKESamxPAgZ1B/FT+18l59DazsMcDXs2/FNBw0rTb31oTgU0gm6rbaybzbFiaGs26k4A
L3BOdPsm8VqblzFbog746wTyTSB/MCFDUuNXJb9bNF46Ls7Xnfwse10wVr23j04di/Bft3mHW5LJ
yQot7XUL9Yk9t/ghgcipon27LOfrgd1fg8sPjzCuyCNgxTEHzRPZid22PGY/02qZyZFsk55vQ/Z0
89o6P/G+oCDif4j6+BDuKxPlYM4OLDHYjQobi63JD94shSrfGsUUHA3aDneUpSb7QmnD88oK3eT+
5eiDSmsIaJ6uZ+Py13HKE/RCeR3NwIljyRoYPCxleFZZ8kUUH/nHHyAGVSCAhYLcHq1qYCPRDH3e
iXlJ/zDdwijoAOpdN1w7tF6TTWbtjPlS9kF5gZyiCtnmmNcbvcEZSyAADaA9mNFMaYTufqmQnQ71
8lMeSx7E7JELDzzQdltmXacSjXwPwxgF+qci5CgToEheVkbltI8n4GkaTC1XiP9vIPtry06TKdr+
1zvrV/zuPALmhF6AoiyyNd0TdWYKahujmToa5EqUYO4elAH9WGEYViv/XhVL0HujT5l4LhnQCYeF
Qs0E93X/0ykQoJPCioyGJbRAilyFONgfET7Ng8Psd/JAYYMGpDkSbMy61gVjwIGUEIXrwSC2defc
fklYTQXf7ysP01kqfsk1hauUAFqgNTk9aCwQTfKxXyfps4qstVVwpUmnS8yBXo6tVD/MmjNVKQvj
BEyP7SL+3W0nCe1RfsR8loiitpRmfvdqY7S6NyQ4RGCf2n9+E+RC64fFp7ybl6tgwUZ8CS6tTGxv
anYmSqMQDUs3s2uvm5Jg+XjMTv87qoVPQtrivgVHnuGeYJkCLQdjdigGJH0FEVz19WQNMeL7oIRh
ErcJ+u2igLaNnUngUHSKFWxzJAY6b3cpKK7IcaQez6d7CfuAbSRQUn4GJKQRG28Gzgh3Tfr/MV8j
UA/LsdZ6NaDvvzzrPdsqNaowXe3id1zUsG+QtuXRj82UyiRd0XUroOX1axqkDtLzumj3NlOcoSd8
5sDbFQL2ujeNtoWETv4uzh+b4bHh595k2sgGwkcXMNFibda/sQwGZ8+YXpIht7N4o9ezG8O1ir8l
Z86mqMZsLU/DoQmhZ+9HzNH2j/k5leemG1oo92gxCfwmU4LAw3rSdPrxbfnKF/N9TJR1khLLie94
g681ZgKN/ALbESMPLU58Z0uhX4OOZTQD/kbqVt0kjy5MklG/ohkfMtmzuD3gQ4yyxX7a4J4asBio
U8LmaRZc6ADJFTTP4fsK/VZvEXDwuq7gpR6DZ3UMVLS9QfTnqK+hKEj4II9eD0uur3fXnsfTcina
DXG8Rexu0pEXUbTVfpbT+qFrhYUewaG8wkuKqjYGOObX0pKkrGg0wyfc5i9PxQmdhZkyBCxOTFoH
Osowxq8gEy0+bnbawlzWUuAOrIbMrZiGIcmTbekIvsgB/nXWx++YrHkusClWqLq6gGpS8y9SMqNf
PfLsfMUSmUkhokHFoLkq12AjnYQEoj51kNAgBOPrNsQZ8dwefLWwhEWqBgQEHGE9VwNISaK+zlfU
5LqyLTkHY8z9uxqknifHOpsLFp6MoDBLyXt6lW6jqNVpFwcFi5yDiHogCnt7K5eIPgQiMMWbxVPt
ykHF1+SiZbaxedq2X4FrbGWHVvV+Dru6e7VvKqEchWCORv52890WKjNmypsoShyl1ac3XOUswsyF
kog/w5cEfvnCeXYshEuFKR3HAvhrpqf1PJgopUZH7582o0+CAvJP28Enil7jrK41uRxC7q2o+oUC
mYL5rRsD4kHZvhc5Wme+74B4tdWK0WXWYdpLMQXOtppbypbxp4Xt2f3KrigBfq7SPRxqhL4o9PRL
HbIofy9QQ0Ym6YVGmcGP5kferCnDXoEotjXgQZzeElscideFc4yO0Bj93L9SmCCERLXP/BwW/qEN
R8O8NkywNQj6G6uh7pgMww3FRTQ+0w7Tngr5yvHN7j7rLRmhn5hXWDWrIDAdiWfNqcNH4OjUWq1o
qCd5R9iI171oKZ8/t6NIhbRoVmvhj9tRxom0d01RxVnN7oqLaehsIkzSdx1LrURyID2EwvMxAD+r
/lTJ+dfpZ3Ybh4EYrssHUveqTflFC5lCPLFtLNqINB7nBkuHYXouuNPowlFNIEzR+AOynKU9iHFW
r6CnD6uLZe0KK+NKZkxwGcctE9kuCgctBC17Ibt7TIsTYTvK7UV8oepDD4MN5Ixbqiba+rlhFSz6
EIimSysl68FXNEuUroZD0r9Q5I3aT77ouF8/OhR0oZhXfZS9rXsPpW2wK/bfH3Chd+BWzUXQkAPP
0shFNelXjP2nSzM+9GitWmGCRun3DFbwOEAB4aB/WtGm36I7pLTqDPCJFH93wpUsMWuU2UGjLR4B
r0UUvnMH8V5GnsyB1ed2s46unbkwVZoGBJWsHdLHF7QddxP6vjiBLsO5sNX5/CFH7yk0B7QRkO8c
x2PNFTYgLUu2qgu75XHU2y5FRTAdcoYH0TdESazsytdiBhDbDBb20YY4u92xQIXamyiGB0tlCv8o
To2oCVbooZWBRO/hVaAaznQ5pjxi0cnZe4YnrBjGDX9YLgBZE9o/zdQBVrvyflobPGB9dmR3DD5K
bSSOu14JS4j9hs9d4lQ30DQ39lha7GAd26Yqq+tgoNFnWacUOPl6BrJy2BTY8G66BZsaIuXdFKrv
eJI9ybI0R4/KdQ9aiCyLG4okFJpKTvYNjpTZm6eJjseiCkpmztbmE682MzXyoFsLnAWD6c64WUSv
y9BSvFcC0eZl7CuLi8GfekTf8hTe8vh9EX2BWwoZMWyB1mvu60pWi29t4P2dHazl6XyC+EXUpBKG
ak7TIC4GR0rsrZ0RNlumqVXbX/rOkeT6I5xoh8iH5jRaNJoe30vrxL0hMyGaW7j362R7i9eGIwFO
/eqh2gZCadYCYzbAi+PkIClq0IyqG+yoIxGulL/7BAOmQNMXE3GIq7VzQNmDmnKcnx01lnkJmmFE
gW2KpUO4RWFvnbYrdnLschl6mzdCp+T/pODoSVfjRGg97gnR4Va55VtwFL/KAVJvwsESx2E8jAhm
IMaELm38Reb6TYIQLnRyI7agzAZQGgRp8Ae++bSqpRFp9wytsxWWJg0LKh4v9FHC/O8anIHqVGt/
GrkdT1WwKOBnFaAto+r0axWwvdIqFk2PYPAzhSEmM8G97aEVJfAkEE6ilBpfbnvuC0Txg93Wr1Dr
4QMF5CvfCgWKICxmhpac5jyWLQDXh/kQbA6xXm9bPYNYDvxbB+Y8YhJ48SBF2HeuMwlkHLvL3OSl
PZjlmQhJcXCgGNKQ7k60Jk3o5Lr4lurjOXyx9mFdLJ83Fy+if4hi+2MfQe0WhcoVW8W5EAtdV5IL
ZKCC2xwgv+vP4HFkJQ19Gdm5t1+Mz0tB5dTYRjowy88yI/eIMx6tnKEc0JX4EBMNUdbauFrXqoeD
Hy887oAu1FueNRib+xPzIWgED42n75bArNXdGz5L3+5mJbQKTPkkfobq0IXdaheCAwM0npQkaut/
fX87L7b5XFIw44rNxAghhxXHk9aMKVClyebNrRl9Bf8IB4/gVsqn6pj+ReIK5wGHwM7UhfkrVdhO
6T+wlkyr7tGlTgdGl//bCTsOswbkUEqsKDfeYiYQqsltm9gCoKJ6O+36g8CVi3D3o4B4hqCHDgTT
XR8jWxw2zszgq9tGoBNZLwV5lQOXnBGTB8UDshe3poTL/3gKXcHTxVhhxIfQLfbHjRmlM08MaYcH
9fSCzvxPXEjsk5SiG+4pK2FQYA87JyFYNhIqaGTSSz1/wEaR0HraqA3du6bbnvjGTJNN2FdA59UI
acEvRPhAv0ha8jIikQGUVv/1Fgiw3/PsA9UUwmc1SjiAfvlAOF+H8vj4pj3K7AiLriCcA3UqLVyM
GozkQBHoVW3ghPkgjgjHxIvTIBXrOaftEZv3/26Oxv9rKoQ0hOmojoxdAYdrt+1w4BkI1Jtyb7su
rB4WeQgYLaKpOKiSC5PWjF0xrMe9t1dTbvSLF4Aztv2m8Lg4znNMTwcifCGWfftuykyKF8sNsyQp
XiIg7mlQHM2gAEVpt21dUVzk6XLGtvHI2NbTNejntscvODcBXW5QMeKVfxsBSgQ0hg2knp6rLekL
S/uL7FeRG1gc5Hr3gG16TlpJOVOnz9myjAYIWkvm6l8AuLglQAx4+vudSQs7AzkHhNc4fTmFXDba
C2goNbQT9qUIBRfmXVqTsNZJq0MapHEZRwQlvr/dPluG81RBf/o7gwvERQ5CyB0xzhqfx+rAycyK
vnR/4UTxO4zT6AamrTn118/t6+tx581bJA5TVPwoMROsYHO+X67WDLyEh08SIuBOnFShyC9NkbZp
RhZc/F9LRqAC0e8RvDFHThyF/HmjHeDtQ95ZO/EUX8JpYieb7DUimHNQ7vLb+ralszvZVKB0yyfg
Ol+LYSgyCUi7hAkJa40bu3S592X8MRciHCJ6U+0HRlWiezd2iTniAZiK7bQ0yZklXdPd8T6ClDI0
U3Bf6B671WPL1+jOc4sN9aQoj+fvAYLKh2O1YYZY7qXM3h2zROkobQ/ONCW3huvHVdM/320PI6jV
5mPIDj8x0JfXUy+b3psMv8WxwPuZxJSOogaJZCOBcf2tyhK2FvKAvLwcDXC/wzVrTeFW9Xzgo9+i
USpZxdiG0gaabWVIKUReuLSGgwXIMKt1v8zfm6awyR8czjkEvKccNs/Ra+X7TSXXoY5FnMIKR7F0
dXK7n0h0Mvd0AyHJMNDK59PSxk5MZqCyy0EFv1Anyc8i1ot/+IVmTJQlepbRjA3w7Yz5W0hpja6F
PFp+Hr3LWFwytM1dOWuQTiLWVKIwas1sSbmVtEsyCN5r8B1iirWjf9lm3qkpsQn8EfkjGypBt03h
bUythCUnO1/g+lP3Pj3dzb0CuP3jZGBGB+Ysld/elai8nDcKBSIlXZUqMiwPaXtsyhGv11RhqWfA
gPJTIRfyOpjAfak5721s2CB2h7B+gm1UX+QQ9YB7YbMNJ0yV8yJO5d7tQycrPX3VTdhpFw3wbbx5
QvGhMRJbSukeauf3JaU0qa/UgAytWHeo2TeeSj154O21Xgk4biWwxh2s6KjhzPmMAfN6/DCeqx0Z
SLY+0yG2uR80QzGxfmXWEHmu0WrBRwx9A5MHC/Bm66dYNnNKZtW4H8cn8J4cEWb+MhD/T4mPQCRv
/gXfN5nOkXu6BXdi98CaJrNvvXkBxmPCkeGvkM7b3aOChwTjB0pI1zqkLj/i4WCs4LTutfbDCrqf
DPLnYoJLqtS92UQISnivRBzLtcWj3u2dmcm5+etXVomk0PdJe0nAP1rnzlAJ0RHOlDYDtU5EKkQp
BB4VWgG6qgo7Zdfh3ARdoL4Sn5NKKlON+xKn+mCpE3ar8ltvNrQpy4U2YuI5CPp9exHs3TYcufFH
Kq1dpL4KM9PxJlMNPA44irGjkyPRdKtdinEP3YnKfLJUfppTYKAuCtViLRf5UrfJ4unX4caUPQ4S
vL1wJQHBZKPmiLD9d668Y1iLNpI7VOzV0uRfAdeXC2+U0yu0eikRNXFSAlMT0vr61Qsy5OKtYdAP
jgxtP5rLz+2MGak1A04Uz/X9+GdgyCBBqGYe9PRWRzMm2FAPue567K/ZD+xXpMF2henCppSfPnpu
XwLH+4xIDtXiF4J05xLa7MN50jhIF1h1EfKlKu3wyaNVJiLS5kexuvq23x0TmhS22a3M2rN5e76g
BA7g8EPa0zhOZjqT7udmEfZuFRGXX0Dfmbdxlwt/OcAAWcQ/H6l6PIy/Q1cC1xq/GYtvGwRjR5GG
Pcd0xfJxxdA/YhE6CU/c671d+wlD10ouZTKpf7SlmEI2tEVqYBF3rG/itG+BjnwCp2sWBAac6WE5
kkWhulmmIVbFHap9qkmxYFll75gjauH67mkgfYvoprSMKDTF0/K4djWdHgHZUoCnvYcjz/uDYCSa
unFqwgCebkMXIwZxgTfVt3LkaZnIG5Jl229QasSzH47qnAzUcBh/cLAKjUbpr2nY6T5MvwRa95iG
x9yssuvSPNB4spnU4uS9pX6OepzHhgiWksNDehXT4M7+lfsFuIVWepIoJepRkswlGWhH8yWrCCtY
rSH8JvOKfKTD8FVq3WZOaXMHtVSW2H11b7ttKiDBCcvrhhzP3cB0othx8OXaWmJpHblA2Doy7Zpl
L6c4xEDvIwObBAPIaek15LLg9+JHEq2kGJ0rHuiCQKjsGlHzVi5QnWF4dRPnla+Aafkwi/jPhZxe
pzrByheAXEj+opEgPbWl2SNIX26P6kvFfNCAv4Dm3vG/Kobsa/NxGltFtIsvY/H5E7JPHLftNFVV
8sBmGT2jQU78hfEJONWyT9efhx2LHGodiiBhRQ2qNQbhFGCo83JkPc/iLaM5u2pbQM3nFvUQR8KG
zLRvhqvvcdeVmAmg8rxUNetkHQW5zbwdZrxgveu0ADar8qtgx5S7EYBaCxKRUsTf48iOEivufI5b
x+SOsFymrn7vu72I28DOfuIEoird82OAH2Hp/fja8038j0WAgNdwGIroz2PzzoqtjoaAFD1flPTW
3hY8ot3WrjxYAl5gryuLutqsINhVaiw9DWLlsoCXA/bfhNZTcg6FQ9QC8Fk62cSOqhViWvb9aBcs
Lc22U6HUwTKQxlOPRSsj3MQMRzBpUAD/pVOWhydeVZ2G21/9yrHPl60FjLdZ6UFIVuaP/dD0pOay
XvyShsrwmIqXajGbggLRe0EgVjuQJ4N0ffkL83tXR8mRpjFEwtUJN5JC91OXSOW8I4n5SWGcyNkK
TlSjVUZDKJlBojpwtk+g1CVi8ZHdfnE0QUcNU/Ckf45qG2L5Kx4n5C0XCVdBse4b3naDTDVr6i+H
FV9gGha8KD6KJWi1l/S1lM41i7vtR4ENPh5kcratVM1Y8QwzDJcAiVKdh5X31HcScpD/h3YdoS+v
bWlRkRgiPXb3FuS+7/4+FrwHqPcVA6WHGMCm6kumFDRcponTn1Z7/q+QakpEk7G0hC795jEJtBDo
m0UDBQ+fBTKmeY9yH2V2pU5ScpZJPYk8/ZBOChIkCWxcRx5CjmBSIhE1crGLo1mnUGCf6qld32pK
XceMIhEu/o7m0lT7Jdkj8JiW3AHp+H+IUngxv8oqixdceCPXXurSJhwjvisUwJezQ24s9mhkRdDW
CYN6uXr2mo5uiLEARfENMUMQuYN6AtK+zT10P+xBK9cR2mbpx7ZD7jOgkeALIH1k7LwxHt/sVMtL
sflvHx6fUACVedW+W4okEPNch8o8Xy6372rpmZOWRYDT4TQFvi3+G0LjWodhXakmnLzCDyw4JNgR
Kdb/8JKyRZpZyHe+PDT/JbqQLUpeJIahsFfVbRWkO2fXXKsm9Nv1kFdsg9aSHkd7nkfnPCT6Ojzj
QgQrke3cbnXKnQyp98H28COhLTWHwuoxIFoAnu9WtD9hUxClJW0kfPylHLCnpA9uCpCG/vDKzQhp
Y5uRBj0kPwTt7Cdg1WmcsOAZMlQ5VtXzFgLzuprZAZWYvuOXBxmQepDhXEQB+KZfd1LlVM0syA6j
vg2KGwvuym2rJvhGZkUaJ67cv3SS7M45GBsoyHm073V3ssTUfznk3HYrDIfi4AUOmj5poINM0+xz
s7+r0DpXOHDc/fBEkVInFESYJJ27DGMro/jTomgpIdnrxoTT9wR+N/+vSizqITeY+D2H1joGxRSX
7uhI0b8izj+2PupyUSmemVrcKCtBKA6/pPUZe4egFS5UOHy1GaNc7WT9mjooYpJXDJlivkW+pTh3
5NbGc6R9zNMaAqpM5ZuYXByFETrA2HvW/LGe7+ugRVFA9zpGRIuhCfvDnI3bW3yPrCDOQSshPaYF
tthKAkRsE8YuwO803i7AgcoXYEmLhUbJruc8BQa6Bj/uu95FFPQnKdFht0V39aaiREUbxlSa0kXp
jvZoGPFH9V0lv9RT1HG7/X1wy9Q77J/F2YaE/Cm/ImQAveCf7fDjWnwuin4Yr1mLByoISVyxZ1wp
TdnPD664lcqIfyzjlnmzTs4aYvCGVJUHr60HaTAHpM9ESEeyr+OdLgmsUNx6/Fu9LGly8Xpjs6Ql
0tulmW4IY9TSdPpikKkkRzKiHfJXcu57DirljfI8I3XqNmK9J67mHEIhFGoK/z1uFJXQxQnnFCpI
uj1cOUqo4LD74CnYvKtKpzWMv8QkzfI7Mkm0NO5UHevDkGcyIE7L+GsST83d+BwOiEjDpmoPN/62
+kpVQKVYCY+ILGGZBO+RVKZojBvMNp/kXUJdABwV+wY0W/MayJNLuz9AY4byOSyDLi715cWwAarg
iKckXKTG3Ot5Cc1H6Vq9wRcQWECKC7Vsl43vTmrpHYYkeSHbV5F9WxzSp+vHOqbOnRqVp0MJiinZ
PONeGp1Cg91aOwXTNUrZCXYSy+zzoACQ3lNPerl+g/FwXwRWCN/QO5nK+KwRhipXIB6oZ2DdaBXn
245UsnrtZihWMIxx24DyEHl8JttLxeIJnBUUhQEONflylSNCTK6eXKb05A/pynjXKERoiM0IobZ4
2bPC5vs7kVYGFpLAMXN4bvDdWs5pfwojDL58vSpZwVYjNt4d0/+/3+6Z9w7NYx8bxoG89oJ7qhIP
AhRMwhGHGazivjYAxuwMOAbZzoWxKOBrk4yCZpKdDg7I74pg50sAxx1rZ/hWiptkLja2AGFFdi4L
1JnM9tz3VluGbekUomfYxOlK5MUk3RQaPvdzmsgzciKinxP23+iVqsYb3nSDn+doK+o2vNtEqKFl
acwf8xmqw46wi77eKrpVKsoi7e6WuUt7Lh9lfP9BGk+emXiLdqsYZE0wRwi4WMdwLkQqf53yFRNP
h0yWxe57QmOGq2eOOfBTvlqTSC5kiXYruMEUUr1ZlllWPEGYSS18447R1h6+6QTw5hak5gQXlLdz
xGLoR1/L5cpgBxGwxOMK9XkCc4OiOMrEP9ixtxfiPBSMVUHdsp5fq9/sf7HOjfuAz8rP+33GpfgN
W3dXOiEhY1WHtJjIpWYg6pQfBeXPif20QnKs6f2yNnGhufqcwaf4HOK5RKkdAD8aDXgyUz5EohZ+
S1GCYZxqjNQMfwWTo8Xe3EnRMiCFci8SSpF2IkVEhoXtU0MifCweLlohqEuVRe4vmNWARAgDE+94
Md4ieQ+sMyrrV8egz8qzjCezN2OdZEfmyTG9jIzwhKZ/rZdkIU6FpjtcmoyOX4OEHT+CuAg0+5mL
ePlMgQV4OZtKfeQjWeQHwICl6LKMBBzaWHWRDIm+I81sBt2H6+Dac+dYV+RfAUOfjFFxP/R89BX2
ZbMsUW30NqszOnoYM3ZWjZYRqMqs9ZJ74YusK1X60tNw033cu1xjeY3tXyw7S6nMuHHVA7rENZ0n
OYjEI1hCR/bMu9RNy7cdcq1OguJ3plVnb5no21fg+bBFpTqNJY86lxVzXxtEiSOu5ZNf5qXsJkgf
qUKElzC5TUYvjEyxHHggKAnqLH5NvFoVay0XMDDVnUO0QVfdJf6CfhMjXrePRMRafeoZno2/45dC
rY+M9Te0z362ljYJCLR2R8Qi/LKIYwqQog3bAYf33VcnmxPLNp8yMkAwMS7Hd2i7jC2JYhATpZtH
NleHRyaT8N+GN78624f+QL4EkuYdvwNTQD2XhyDj2H+YVnJIDqayckixV0Rc6UwkHiMGTshbcEP8
A1EiUYjti5k6ylPsKLt5JCwYoaz+/heFZxd6UOUfpGCrmfxOTuG5fFniL+8R+jYZDGtz1sHLktn/
HbYztYCLK35XEYaDYHzncyHRFFvfFq8SGPcOufhMmr94DhaFfpX2YTVAkhz7VBJUxtNdcEkHvzGq
XI5WvpVYsHOiLfg4oe9+mdbXpGAGQmlJx4Wy/g4Muj9+0VY3Z+FQKd64ZtjbWZujmatOY8J0bO4c
uTBHSXXfzb13MgfQnDD7j0Gxos0s/dHuNPAe7rt4+11ok4WokGJjICx7CMIzFls0LBh45o4Kwl0z
0G3BmiNP/CU56u1o3tSMO+7cGXJhxV9wv06RIDtjY+AO4ZWXdpBTcyOVR+S0TmGFImbDvQW8PXyB
kVY/AcY5a4G4ZWIXXuMn4IzpgU6BamWv8u4nozQbl8ejWexSEPJ/zTZnftKhMViIurmsnV2cBBxG
nrb6AhnoC4hGccDHlivStR6dbjJE0gt6tIDRvcStnUSF4QMUS4781LPzHkVoiPuCL0JxN9epB5Pd
lxdcInkEIwiq+ru4NyWf3BN0Y1Ut8NWH4X+Hg25pYBlbj/csHY0O0OKroePVnlOMWQRLaOB9WvBN
xhJf1BRc+2EVX3WzMSPdCN39BrUXNlZEXpwMkpmGiZisVpncvG+urG8/Nzw0bYAswmtPc7U5Lm1T
IZiLmhrC/9reCM22EsqKl8HH0CHigVruaOz1j4wW9NJm+/ytcuNoMHzYlm4zZGGGDZp2FTNTTnM/
vHn8zDfh7A/l+PA62d3tQ9vfquYWZb3Mc2S7LixypbclJwevBxbUWTZip8Uqp4rcsl037bqpnB0l
IHCi3HX0wlQT5DKSJ0O/J3S0aH0/vqNglyulmyLiU+j1Ckvb+TawVRC52J+S0xpSp/t2uO6iZdDc
DEoFNjIpmY/H3Ge4YJV9QKQ4S2CKcPLBNt70V0J1Ve/WQZVAmdUXluI+ot/cXIwJ+50edw/ksJ4o
+QW3PZkzFmt6O4AoReX3VzW7AmGczsCteu+H038G/ToDTGfyM6+Te3ec6sdMrc1D95G4qA69AqiF
Xuf5dHzeiozuoYmm+1jbsKtIdpmpYGe4Xz55DkaLa5JjV1ZERhuNx6tullKv30YGeTLUtTBi8bGg
2QB3QwFjujsQDBcSywJn4B9p1sQ/gezzBBKQ8q0Qzn6wppzIzgu+MzJrfncAqwGvLXmz+lfpPfk/
fyJe+mbMXztWeLqVz8RLjDIdMQTbq1Pi92cZrRpMYvbSbm7DtaFymprtQrGhAThzhPduGYygSPsI
QPO1Rxv/E/WMLrNGxbgsyKWiViPwakfIRUmOHMPjapS9ygOah6KViuiDAcg4oL3tFCr4JWQeTuax
a9qtRya54OK1OvvksTiD7NHgV0ObMyfEH8aNAPWKlpyzQ+rr9zKE7g+AA5357gtELoaztjFXCEuL
aWWL/qaar1zNzOHo6h9Jt7D1n0lxSZ49tJc0LHztv11hRJQAWECL5Y3Nv8blFdiDJGqtH03pAF9y
TmRSIbNi/IrRTDP2mfPzgX0ZbTTun3cz4o+ByYqUsscco6/BLJlAdCku6mNCf2ft8jXqv9T6LVrN
XrofLH9scWCf40ztAi5u
`protect end_protected
