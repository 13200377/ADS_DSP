-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Y8PZgE//wDaIdA1A2ARqf/qUQbjW+ghT3U/YNp4lcUT87xSkBIEXQLUY0qDduDopXZR4jG8Ba4EV
xGaOjtWeEflzOpfeGgf3vuH9TtZwkZQKbStRKE5dvpNtFru13s0SoaWk2EyO+rkZCETS4U2jA/4Y
WImJPqcaOb7mcwcMk71v7G+/OsuVQkCkBHcKYf0+wzk9Wj89Sl9oozYW2hN7HCTyh5b9GFKvFppJ
mJt/aj0lfXkwqsTY8I3b6b2U4x+p0xB9yadTxozMKs/x6EbChb+gy+ogxAZbzUmP+I3n+0IIHhRf
t205MAngBl8x4fScWZbXossXBTx6ne/nDJfb3A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 17008)
`protect data_block
96fBoYWWTDaCmOvW1kbvL4EjC2XhIL6dhrsVN3BzhKPrpyAETQyuWHJUWhfmS8Gy4zNlg3GFrLnS
mFTirvaWF4meKAOTwqx03062cWkQhfpkTOshW54gOvzK3J1TCvNKIXPSP76mwB5bDYD2GQy9TSHw
VI3RsSVadmULcCqnEungBc5q5fVngguPXBa1Pug/ViCD1xm6pbL8BUyXNv9fQGYW5g76Y/xRbbkX
xFlRcOFrC0EapOwv13Q6anazFbP1qDTai7/Cx3pljMGmQtgCcL7sHVZsvvswjN0WOengQz3rxgPq
h0lvgYtt75ipDMCNvnmntzw6StGS23Yah+MCzaciTcdwEnAZ4jT8t3JPLR8yHs13HLuAhukFU42R
1gxz27YzzwmGbqW5h5Tans4mgQeA/jrLUmGD+0E04ubO9AWVpRGJHMMi6I/UxFw0cjCyhK6LYzZy
nWlZrSFwWI7k369UqpbTIyIb7z6AnDLnLKAOqKehs0ShFllRUhHjAM7rldCNsang0y/h2bYlHAcL
xYPbIo8kiuANAg09+AgRwuD8Hspo/n++rbzROl8XYbld7xK3sFwsyBc8ArIoyNgKiAmw3BoPrsMp
AoUAm5IWnRuthv/NVS3ZR45mKtuJ6iZHu0aTC0eZLMHvpM8J6Tkd8leXE932XYaPydeej7BJxvop
AIjWFLHKGpBrwtTO2MkspPkYZCXDfignLPcD2GWvArRa7+qXt42k8dpHpy3Xc5KgpneigkQwKFBo
5lP/tfLNb1BDRuE90g4T+GZy1QXPyfqTqmZiTxjebdHxGB9TGYXBFXugOjSf+No56IvbjNXIA42Z
d3ol65ea/pB8yWsO34me+vbtSbOW/rmuTpeQdAYZKVBWUfevqYqRcGtkOLY8MJlTfobUGTwv0T/W
Ilgb8bF+yVPq629XjFfAoChrQZrjRw9DMg+4xQ2zXQAIat9MGVNsC7ejDKHCtc2tM5qYbJraI/LM
C45C/a96B408OTXfgldaa7Pq1BU4RuAAHtanUO/1a+DxXYl8l2GRdq1v5ACQtoWgnDq9vdFwBglm
oG4NQfYn/eQI2kxLX9ESy2oGbj9qk9ZunAHuRTjDuewb4n9+G9PCUlCHIZxngSMG1AuHQgJal/Pp
OiGcIXU+17v1NguTCib88/iL5HNa6Qko+qGs8k/DwfIHQXZ96cumTXNcYFjUvi3ksspSNFeZ+tUo
23KC+o9NB646kKKFepFcsvwfganrYnmg2zwsMnHWt1jfspglG811YIvrABKf66pX53s0w4u/aOYl
o9NyYTxQKQD0Sf8k4IeAssaD2CxZvH2XBcNk58YYP9KLLVAdGCMz7Y0Rw4QoUR9D0skiqPXvzH29
sj+aiQySMzyOdXfw17NN3+TjxfcrP4wnz3DAq6GJJrIBsAP6N7H7WDwzjeIdKg5ffZGpSVIM2Y+A
kXna9F0GpJqEq7o4AggOp5lONPi3Ezj3fzkNjV8DYaMXRHJHh+RJQJUZJKoAJWAa8JpWB6NlpY7y
+0PMXswy7FfzQaLZ+URu8TiCfjSVuYvIUIr+vQPVpCbBALdQj7tUzYxZMffiUhfN6cO6NB9S2gi2
vbuWTvxZMq5FAAQjR9ydREcX3Xn+sQUEo00EFH34P9flRYNl0GQvEaGlQZSeYd9H6kIt6oLbVlY1
UpReGkkFh4fiHUIACtl5ZUVsV20SetDwMbzzotjTFfOLwnfFMcEe0l36oE9S2yVXngaXR2Bo80x4
tjmMQDFHibX55aoxlRk9uOdXLZbKGWBlgNCvxgSXf0gdMDHKNDV8Drw5n9A9q8EPR5c9tQkZ+wEu
J2pvIJSU/SvWl6AuFYVoo8kp8lXZ8UEcxfgNoteXv9HguEoznPrzjntNSCPPqOPraWC9JD1KuSNP
Hna8jzX51G8mYBG9FsuAq+zRDk624LrD+GNm7z5otVfbQ8s76xRWneOQ0dVBxZoYiDkYmGaCZ/tI
KzRqhVKMajwYkO1dQqUXLHzEOitlDhN45fSNgM0j4O8OTaPu+q/6+y3YjrUTAq8nJnG77+xXS2Hx
9r0z88IzhxXHrdbUlY/t5KjES56Q57FF9s5z/SIbCxd6EeFaerYxw4rdsd6wbFnfWSqYZAatwcK5
CLn0x49fVF/f9CYQewxgJ1khwBjvoMitmvpJmjqib5iSn2/JR8VYEcqpArHRRg1p3RGR4i6bimJl
ovtr+OIFOv4o0n7kdP+ceYMAm6kIi7PiKSRxEKEwVRQ/yBe+Jmg10EqLuY/LCGxn9DHKBkXpSOJr
nW4M1MXcovfMwdowzYAJ3Li4jWJB6xaP9kYUExg/ttVYIPkmdJrplsF5Fo9LiCts2GLGxxcI09TP
4JtN8qgtvnE6VRWTgGSzSniB5g3fMDCapWhN7Tfzl/bGuoflWt7Dbw3xZjl8h2QneyIdBOmEqdnS
7WmLp3pc0a+eyQoyfcO/zZCRCwfItV5Mgksrcvu2GuHzJ7APvYiMhWBx+vKMeOdo8lMhZdt557IQ
Y8VZG0H8bsjLL934FNr6NtIrJFwmjImKHzPnmDnzyBRk4sSLxj4QjjvVAJnthDee1YW+bYrdFpNy
v4KP+KxNQqCGNcHUJMOxv7ZI0qrci6tpJMc3yT6wVOvkPryGrj2Ip2m94ydRVczUbwYjW9dIo69/
Mq2wQfSyFSu4SVVmbxsX61VXnESx1zQuX+fI0iK4JR03HGvhmDEpT0mSvCBEXObm6837lvF0HV6P
QepJwPhYk1858RU/QRaIyX4cqqxOBz4bHrVFN85vC0oqpjYfu9QxO/YzJNMwYYHlaG/+nC0idWLa
mTE8flneQqApQSWUub+7WE88iDkXdXdCEWjSEMIhOuF0QhUOFWqV2xLbOOicdbKloTkAVw8erXO3
ue6WhYOZgisDU1T3Jvt+aScyENGKjsDSV6rma+jbyPtrUDj31rKMG4IfaOOO548G5fv7P5QfdSaJ
BCoUGNnLDYV/TJeb5yWxCRc2eyBCE0P/B913cGSQ/E+HOfwXQw/FWLp9cXxcbz2fzuuzguMFUHTu
lAGrhlD9IGYcAiLoXcEG9W8YHZsqqEe2N0yVaw2Ps2/AIOyemK7HwNOP8YwsSAxiE042hZHTgvad
s9HUBLrog0pUxlnlr1rH0kvacdLaUKo6qgBbVlH2q+htXWpubTaZ2ZY9kYpndAszxkyDT61tDgBQ
Q0zH8NtwOzb1I2bcQZpC5VmBJmDVe6O4RWCBXobaiLUn1XZkCnTf/C1tbYkIoDGB1bNu7/HpIsDt
C9N/xi4ozCIQEKYAA5VZ6n+/F04TSKmy0dF2d64wJ/Dk7ksq9e5D9VBok+8NJIAkujemt3sU7HwG
d7nOoVuBQX4v5pA+muqFybacSc45ctNRz282oypOAT5k4PhDaIbCMg6USuMQPhDcn4gtJZmdPsCl
1CHFFsYHR5gX7QbIVanJu/gyihdBx5/+U1YCQbCqNUGBIcaVYJhaLnftAVV5cukuNUWTUssmXKfk
kn2QDsyjYz9k35nqA7m6wqRNr5L2vaIe0GqREMHLN2OhNtIygZFiJ5c0ugvO9uq9AdSqCZZ6ICl6
BZJD4IuNA4CZioz4casAlq/VSi90Qg1neloX+hUngUpDGOH94z7SEVr4n10ddK0cbZfTPjT6ttdf
UPEqnH2/+wFVAh3WYtUnxGk0AVfmShxfVXd0nhG/FOBwsd4jE87xy6kKgsZmPAQf6ud5oIdcpAbL
vtbSQl/Fi6UYFz+arqTMBaSlKeGo+aHi4zA6n6rb0j86Kn8kkwRtLAYezcf/D+ePuWSlWRmfG+1m
OxCiaqn98Y7Jo00syrgNTSl8KMAgLfjGjYYd8oDaaEHAX2toUvX/mWY9mgSowFzMuKusZha5Y0Gt
BBlz1SH3MhlxrEK6JXiaSaW29lIn8rhasT4QXHgBzoTi3JA4R6yEaHfk9CJQBnHe8waiepEuGE93
7dn2FbIQKxgMV9+I+PZKTh87vmgXlHV/utNxL0k3C6q5N94oAOFeiGRm9QzepqnY2U2sRkL2RKgc
vNR1nyzA04ZVRxkYbAvzC5C21hWA9tbU8Ou/M+XFzaFiwnW5yf5a9TDbr0dC6dBEsqcw92PUlOZk
ta5Kvo9Ilg4SJYpDqoUHVcqICyWbFdmJjQycspEqtw5VfpOZD77Yjr8iVd9wic6r5n4kT4ItCleY
Au1Ny/XlQcpakjyGr7MnWg2n6MDcW+Pnr5Avl7x/Sgs4kSVzGyugB8nhLXW3L3peBVRordfiIMbO
tW3VkIGiSi374s17T15Y75n1v964GMnGe/phGWt4X9McfkFyCT2U1GasMJq1Wma6tliUysP63KLB
MdLH/LWqGzHMD7ZQpK5SH36lM6pDj0D2s4oihOBVQZj5BjGkNDwdLM699ALAAEvbCgFj6zu84hXO
PgAQEUCR8SRfEwzkAP4eo/nx1QxmeN0mFw5X1mAYm8QQCe5mqzo2cAdlEFaBn4OOnuLfJjf6OsT7
eDX56cbFZRmSOXuc+qUn6Mh+I6aIz47rtpzs2mX4EvDZ4eRkhri6LyqY1dnzpAP0JabMjBftdUhd
+eoLo8mmAZa5R2gWDG91Yj8y5YMi+Peq0nBP3MWWMubqdaQz2kmmMRRNPS3GQGQbj/cCasERKFVb
q4smIP0E/dKlU+aCO1CiLrLrvZ5lH7HXPScNtJUtb7nxfqeIEZkmAnk1fgOacTe6FV6yg60Somd4
7FI8A3pfwWPSCQZIC5gLyhX72VayCBc0Gq/j5hiqZ0qRgWrdKVOKvXA/fwSfBoRcYL2gSnjGYhcY
uo6HkQzcDngSy5EhdOrQyKkDWxDe8bSaU0eEJUPOc7sBX+GZkzXUqJ9jJK2mpsyDhAxzhN59cifI
WPViJoLRAYO26avAaJj3i/7ondpft91xgtdjPgORxK1b2HlW6NAd3AJR+Nuv4JR4cKC3/k71M8Vk
dW1fPJJjzK4rvslI75RZXkByiHASKHjnShco4MkMgMxxAOP5oS6sJX2xYJVPND7UKO38DRi0ylFl
UbVJ6uZWbZ1+CF/54QEJ+bVSApmLbtuQcHyNkeB//xy0Jj8rtfkIGswLfOFRERwzZw4XIcJsVlDf
wdsSrbHjriK4pCLy88V7UNfqE6OvPUlJwRWD4/wiswI85CLX1wIauQ/yVNHkIu+ZWnGHiXoHqsIh
VFi9vutcmoZT6cHQJFvpRGZ4mPtw4QwXSzO9/j083f+gCRzpXXhr0SaQag1CcFOtZZot6QHJmh10
V3+DHWmDqoAkXhy+MSzzfu1wgYzzSJCrd7YRr2+nme8dWgZKavApG2QKe6wG5NPoxSNuvIhGcNWo
N1Nr3eDthjvbvg51I3GPu+L7yiPXtzF4j29l35G9LsmAodNrCb3cOtgpcaERLKhQaoae2A+XsQqn
Kfq2sxIv3EldRsfuOBTGgGKTBF4vtQnEoFI25FW3W2Uqc6WkpvQXmhX4lQby5gvL1/YyweHz1Q0N
pLDwCr8wBnhbzgziZRpizdwpzlmaTmZeHxacTq//z+wo5SDL6IyWaFCSKZuA2RfS283t8raaR2Mj
5QsyyM50Bfmy21/2xb9ErD3izM/zpd/3eNxGGD82zcWC0l/Oqk873srCgHgI7nC+Z7y4prrnVdoY
I8fwNMkLSSbbLb6Bhb33x5UnQ+CGT/Z6XAhyrc5t90wxiK44KXreXuKZO8RYM/ppmJ+UU9Kspz12
JKyHQDWj4gdXLq2gILCxJBYgBJm8ioibSWnG8fnv86LTkn0UMDVqZuWFQXJ3nnwPCopCbjPiPjAt
P3C05BQVqsGGM01T+98tGIKi0lfGgPEzAGsU/ffYVOd3M0HxJiWlTE7y0tWq06eBZJ49dP2G8zkL
gnlVvIQIB3xGMpCPQ4hIxzp0uxEvh09HV94X6VdCSQlvDjQ6ks36XsuA0MGQIGT3FAR/2asTBZXa
FzHZ2mn9oeXB8lpErrUcItMfxODgdkBhmjy5r0Un6Sx47/wvgLXginDejq1iKzRBGyzNxH9DOp+f
Y2WwX/uvgOrRDW8mO0VQDIXNKkhf0b/eshW2kJ24cKS0g9W976uB24X5j8bOV2owyAgLu+lQ05C7
6J9oa6fgQBJI/KNgIRimPRVUYDi2JY2Z8bmIRJw5lsl0W/JNoVyRhsUjfxoOBuOZFxINURnT4o9x
3/qIcujgOZXi1c9fNK/T5xGK/kBzVCShR2KXxlkKd5aenEUTUJCw4LzmwMBmkYuIY+4l+iEmbLnI
rXwvcRu9vImi7rLvvnoXUMMCM4Y43APnhcvIU6wURO06y+18vxYPROPoPsaw8MB2t0Y+uSL1RfkX
1glax7ziCQvq4Fjy7Brc/MzJ4IGZYr7n8Uo5MkRJb0uPqMrncZYYZYfz4a9F1MjOsANZ/mOMb+dR
laS2UWUsUe1TxxSH2dzZMLzl/tWw13lxLVpnmrWlQaJO5Q5ssx1EtKm/pCkoCr3/ykHaizAifvPh
goBIf/jYTKuSrOu13WFgtAUJJuuAwHoAzac6795zPe+RIL0JLIvk76KGNDHVfzLUhfv9Ro6DdEF6
Jl8tcNbpHSSjrL7R0226pV1q58Q+bGE+2Sc3Ufh72TQzqkILyGDPZ4Fzl0frANV81FOIRgkGCiWC
g4YmfiVA5Rk8/uOW+tqqvU3R/s/ZFDGUR4eMJLTS3Kruy0qV34l7oJXrW9rKPqvuL1dWha994ckZ
RrYIOfSuOVqOPJCxBLw5unu+msyJ5FB5UIIzAxgE+pRDrJj1epj3zdtq3X4rUr8+PD0LRbFzYd9t
V4FaiVqe+t+0efSaJHXHC+mB0elZ1yMRhAlkFgoWciXfm5FMrkhvCp5oGLThmrMZm/rOJTGuoLzj
AheKOjZqqE4dBdDjG2J3k8FQJf2iBSO8Mtwb2Uj9I8B9MmOrY8QR+n/acMDA4MQ85X6QzBUOojxU
sEyqXckNMX6wKojNlE8z93xCNq3EhWMr9aIpK7lBQiUWIOtZX05VPSHxvZ6t5u40fNJckK74E3UC
k4x4eYYhSavX4Dpa1o+syWhloMgxWQZVYyP2jwAD2ve3uNohPDjMA+5xT5/Ip6SUEiWpFIyO5POd
8pCa7GbAKwDIqlGVZz3p1DJWMl4bbUcV01Dw1M5U0aKrwW7wQzacFHvvttWZBKuczxlY7YZ8erhK
YXjlw+m0JdC4Ni8BpjKHlMpr9wGS8n1fvL/OfzWTWAFVVvM7/NEDcBIRUyi1vcc/SqMyBGWpiXne
hhqi9/x+8nFwnBwSoXSkWN2ShYiU56wV5Qs7SKO4l4ZME3wwD8TYD16j7HI/rNOFf0e4cO+AIlvD
5W/fsrZYO7BqAKR+DGs0JZ/RP6JWIDP4tPsQGlwGnc3+HbY7atuCm6uB61r1laoLd5eoTiv7B9PW
4vvhlz8uSl7DuNiRzE97ZYPJFSFTDxrY6ishNOgU6h1N/ERYm0icxecWlQw4Sqx4rMPABkxC8diH
C+/K29jD0xQeHEiW86et8g3ewUD0rB6S1PCYTixJBdi0HzlMEcmL+o8B3Kmon4459evXyGYThqNk
O+LwImre02fKW93Ay3S6PnEjWdOJkk7govHqEtqfcMk4kHlAxMc/MQpUYPoOGx3y2h5FSqL4sYNx
Q+hvPeTrNI66SOkFt6G9Q72+Nf6uBWdFSpI5bX5TK2dVQBOX+zfpJBIRRbu7rZz7TUemiZkDO7pt
HYmDs6axnEMBhts8swTao0kLteQKvXnTBq7xTn0S789T9ZhgTIKTXs2Aub2shfs3tXzhwwSxk5hu
rz0VHQLYshJ6nhh4CuS0eJ3K9OGffuw37g3k9Kk7QWQImEObByLPOem4tNaxGhxS1g66VYV/gZt1
RVOU1bSI2914qWIwV5YRwC/ev3kNRZa3Cw9yz4mbQqdXahxSVnzxZlUKDSyYaKs037nNUna8JtIG
mbQ1H/WHCLRzCFgzmypOGRcZ+nYI0L2Z1Ric07TWzIdjdB22yd8sIHPHKx/tCJVdz4VDTQAjHAWs
GsSi0YUaVvMdDM87GKFoLx16ACecpywAtJyNu3R+uepmxuBtKbjlRR44TlKTeI/IMaKukU991eQe
lQ1o+NoJSDXx89dXfKJuqdgrPtlYmS3vGHyOYzMfnphr9M01dkt6s6aIB5AG8Bo1vV7aQWa+JNOw
RuxJj0PyMzf9+ZZfthBIeuQH2HEpOnIYLe1mhU+06bZOME1zjCzmbF2qrachX5T6pBmjLCnRkqqY
R7v/FTgfep/i/T66aers0/Akr5UlUJrq9SGdvxbgv/HlFhEwMIWCb3ctVDzk8bPb8VY/2XNZEraG
1F25pMO2WbLz9Lu+T9BWzmdgjQzVWZ6wD/tREPUzcYhuhk1JPvsylj5eJm+l66XkRAnSJVOTnqsB
gV3q3eWX3BoE/pDdNy4gqz0YuhWZppw8WBH/IlRtUkuidObrAz2BMPw1NWzRME5PeDAjyLlz23mr
U0ZM6LR1T0sTBl+k0EpGhr0JJWEP3xMaWxnRnYOh2V69pVOWUe6mGefAhxbsVK8d8Gmc752LkMRb
jpfOp8+WAV6PBaH9Ce9wz/zKhvWWP1gflHUYj3p1tq+bE47r8hqc2/8K2QVVwYSbvfPw0+jUh6hK
GDyPYvsAoAmQiuskx+8st/EBrze2uSSNYhfHBVipxW+2MK0psZSkQOPAYJiPZGaW75Sc9u2IRhj9
psT28UK5mXPqRdnqSpo138LBeczZWZD7Eoo25Yr3sNR96fTttjhNn2h6YTr3cqC9Sgm/s8maXWAl
cs7O1lUkHGLoOgxxoRdxhKBkf80DhrnSU1rFG2bM2joPN/2my1kkfu57Alq5j5OUjm9/cabkS0AU
gd1+l61NQAy/UKWt7g4DhDu8K44sawmNuDU9qA2N7dDR7TBF+BVjOwN4ozN7hQJyppZotgmQe3jn
0B0kEs37d74MXkNMJoyI0+PGGS6nUXTkqQZYh1LjVdy76SHD/wqnMQKxXLLDtWqrX/XE57IGiHCb
yBrj4HBtmeUhMV+PINGNCB1KwbbDaXVyssdFVmivhkz2WsIk0sYCwswHCQau8mmUpazRin73Easp
6VONYARBdE103wga8LajQX80HZHpxjZ2Qsu5lFTssLpUbCmyu2QcAhB04quB2wCXG4qAHq3L9GdV
3m7qcWP1p4Y5Q7sQ0vAFeDSzjwK1JY5CWNsdlWDm82wvBTYQXhvH9BMbyhzmxJzcodHM3QEUDAus
Op9/NyWjh7Wkvk4v7d5Fciuv0KF9hJtZQSvTbnM43EL6RxBq7vmd8vJj9/x7CaxyQFxJwS8hB7ap
E7aSyiHhmu80lpyI624uOip7hKdQanyv97D7pEANj2AFCpfJWDiceMYd/OU8FXmCMNKxzxAZPkgZ
IYsuDOrcc1M+fKadOuovAOVwoEae64Of8MaPua2rdgL67znufGkKxRhUwnJC0EFLiKIvIzBIBhFU
jTpby3b1uqhNywuAgB4nUHpq0APjE1CRYUcpWzpfMN8glTmapSPyMtecZjiUwMB6VooqgFXrYp1m
Jg2Ch3Xqbtyp70pWGxaC+tG4lpOQ97+AI2obVmwXLv3J0ctXA13gcLOf7ffG0wSicmwKsgd13Ode
bHQFpk58Vr9K5O1JwuAym4eob1PT7g5zH84xtoa5eB/QLExIb3mg4TkCe9y2oUIeaosFRlDAvr6n
TzPhHJF2lxGJdajelSpOcfaeywJ7omMu2zOaFt3HBENWBpsalve6l/7CyraM0yT07ZMGT084dhmR
M+sd1VxvPQcioWYqfVVqv2A4IFWvSAxLp7GxFw1dxcPtea7qXg8DkZ4A3/yXf/Ku2RU75CQxrZo+
Qefn0CMeSJjH7hE8xwlojsxg994GRHj2a4vavqhZz+ocTgtaZO3ermngXKzS2Jwizr3UEY8zZlEH
3T+gc+786d0lgJPqA0Eea6xLLa5cVlEX57XB9agiQbH7DnvQdW3cJYVIU8H2TbQjFF/AIBA3AaA/
rpa+jU62BtspMp5LkCN9dAwSFYwzvDLRZfpYWhBoOg7dOaUGKwTFV0Qg5+lguTEP3Q9TqhdLTQHp
YYGw4ATTMc/hVhNUtZuPW1N/dk2zQ/gxg+5OJq9A+Y2+VhF4zuXSrTrj8I3Zs44jRf3Ze7CCnnWq
P7+Axq3Y578REpuYrpLcVZqYNpoTUk+LV4clVGHE+apEcDVmFjSZdujiWRlWzvRAqwlfhs6q+unO
esNaeuNaEjvjuE/xalTrK+psw3/aqYV7jpS7QY7bFJo1tUNjwcKjIXOemaw/b0Ksz3z0Cdn174Hs
PW7W8xL5sZfuUd/Bor4jVf/dOdc8PjKHosDUG6F/wq5UDE0QgdVszjLziJpT2VMEgXDe7AGIMib1
aR0Yj2n7eCi0PlvsIlRNLSbDGyPZw1+RZrNWZVEbVhoH1EmT5uwpvRWI+mPChafvAXyprHuEp8FC
V7pkwqfqS+gIisNfars2HN2d3LiD3rh9MOvJNsRqQEwJIlKXKc/K3kTRFMLbegWiN/iZ0YXD7Wyi
R0/jvF6T9WzlKrDi7pKn0jqqxfNMBFMO7h8Azoqn11JgfQhOjpSSbBIhV04fDSgvG4h6f4n4Eb5H
eAJVoQz34DqAYnvZbweEPLWX4TL0S/NwXHSHOkpw72Vw/ePnbZkwfxsB1eIFu0SZ6hx5sl9TPoBI
EropVU7ivfPDc0Oe9vfMgBPbiO9gfKDYqb4uSjzj08AbNgphLfaeMVEvXFcX5KPBYo9KkTz0H28K
uaSskzSiOHm8oEI592hIqf0eMxF015UbcXD27ZPnjJF03i2Gauu7qZUki0+C3KKD4fjxUTOn8mX5
kilYbYbBj/QjYBIDGSwKs6sh7byQotlkjW36vQzX64VzdOC1o+DsRRQXgZJJu+3qLe7PKry7qXn+
pyafscfm3zPbrbj/pifYASeEVrDdtf8mCbEp9QKx8/xyCRpH1Um+VJCwAelx3VqrE8ZSSzbvl91a
npQnbQWj+S/n9dFzw9NN7/uRnWxRr7POhQz/JIPnzmmfmTNqaX4hOsfSiKxGokLB3bPUKpIDWOIx
33QNK4VYCLNjH1Vce6OOt9hKZdeWDqRO2oevDWDLEWnfq5hg/ta7B5STfjQxQGXwOjUtI/Jf79Yt
4RU9GzIDFP1LbXisPniWtALvUNmkAeVpGvECIGCw5L0MGrRaeGlMy5fJh8bhUScYPsYJq8nacyrF
7eDXHd5/1Eb6ChArmcsNQ/I7Tx20mBe7JeWPEoSbwyMUxJkfHftvZ+kM3ZqegKGanJql2LchB/6o
/z5U5m31kg4xFxB/HsMH4VgryNZkdHNAn1wqKd6iKslCIzncLm/m1bd9FC6W0Kyz2qsqP6o4hjUT
EzEbyQqrBCnme+ErqfETKAy/012+w2DEA0gITxPhzv3hZPjrxONoQe6C9xoXuTRYSSWu3owgewBd
ikVb/WYMMlkQTEJJoydS2yhibN3eWQ5roKRIDlrEh7zGmoI4clywuSz5EL01YbcwMZ+EzCmm1b/Q
RL94q6OcE00bXHYEv8RXs8vHeKU2XehACJJxUxZRCn8gJexH0bPn4Ozlwictf67wG3q/Zd4nxZuJ
881ut+0W+RAziJgvSaSiSqFNq+RkfT9KdAYojqBm/JZWoleufbUPDIFhaMW38rTGS21OMpq+XJoZ
SuUpNwQfIKdHZN1+FqzX/asD40Z6cDy5lKT3sbTOJKNP1x69HuvZzxsqV/0kP76X76KKyC8Vhfde
8cqfOwXg5r7f5BzA61a9DajtEoJSEIBXttXw3u2KC6xwwX4rpGidfYVScYg+Z/JNlmwd7g4mCL5o
+W8TkeXYrDTx16prFzVdzjYIcygoiPsDN7KJNGkFUXWs20HCwIb1ScpKNKxHhX5pUeaWgHA9fS3U
qkXaZz9n/5KdmO8xH2pBMhrzp/ENGJYQ1cflBdBRTestHpAUCyvBbDi2eSQiQhl9ltJqd0Q/Hz3S
saJB8r7iba7hcbHZDxqL5pMu8um6R4fpZ3rmzVnVybMRkt0vXJrLLoopQUgj0/8gOhBENbh2TI4O
qxR0gtvMRTRTCfuCZDGQPVSBN+2u27dp/GTYJPgq/0LrLrg2l5sIeZ/84JvKDQU2wrKFgeN6Qd1F
hHa43DAPQ/sWvE2cxAw3r8ybgN+nEK9G+qci/4s83eVC4t7LwtopTAsO8CzzBksfRQS8HbNkUOVI
kXis9vAUdN9lUzXwimOBaOytpNOaJBW34xDfSoqelTl69YFtNyaVJ6fNq6j7TRzcqWsXLFqJbom4
0hWWKlxaO3YHu3bTTadnCsnV9qfBWyh9BCgtsXGWGC9f2UVVgJimdCSI6BNwuFEO80WBx8lCUfeq
4zdDBeLx8s/2j0Rt4BXTFxaoMeUVhltwLnLY9PphEv5hoNy4JVba0VBWMFf/29TgST4DtN29FEtm
HYfrYuPsatWjkB+k2EHq02mgbzTml988lyq6DZoQromLya0LSqPwPeb6kbgan440yl4Z7TlO8xpc
jqHM/qjfLwwwwMkZoGQ5Ca6lXaeOOT27jKw0CukRihDDTQmY2+YE5UU73q8rHcU5nQ8/QRsql461
+z6PRj1rWhNtXBuEY9vjLfTpVfxieHY3wHF6pOzmLOeVZV5WwhWf4pJi7hZO0Soe8DYrl3W7cM9z
VBzAWuGpNCTukIr/IGAaFIHyzHhUtsTxSbxvw+Z2ON2hQNJSHKsn2DK5hNgGD4GXwVktq1myZSvU
NpRxtRRQmhfFLOMNrMQ32pJYgawTnc2h36FxTG8AYSdoLl0B43y9byCR0Mru2teyE3S0GtCjRkq1
6VMUhv0fGoTa6EHK3aGypYP1U1Q2FGQ41ix66r7NN0pSGSZ3X2qSxSBHjiFkBpZGFz2AzN/nMUvN
hDT3GIjDJb0EerVXGb96TjAqwOrTxKAr/Q3JY43ZfEMMTWmxnZzl5kVQ2dxaJbpgtTW7mLvkevFB
IxVgasBI6KWyH/xtmbMNLb2kTPDMmxIicN+6+LFB1HNkxUY+Rt+X4XF4xmantBoFjDR0FToOD9s7
VxLGWjA8t6cTfGrjVmssaZibZIKbq2oBgL7xz2Seu/jJh2IBvDdIxa1PF5hcY9q4Adb1klSFgY8r
Qrw6xgq8ALXCT+6xWXPZ5bG7NTMGfMn06GVlsOJ6pBWqWd9fVFj7boBwAGP9ru3qK8g4GonPdZji
uPx/tViIMHZHWaKbP6FjfuNvW2bsGqD3vUy1jB1VRFUUrVeevJjNia+67NS1sGYEnJ27vQF+VhUb
1PfwSbkU0ZG2Lr9Oe17weWeRwUVqGdX3TNx8AduJfUlRii+78WYCWA/M1vzX/UPbbHNv2Srj1TNN
OYrkncj5Tayn2EGOAZF9+Ki2qmEENMqL1OVmojG84tj+Icwyl2d/LP5kw1iEKfbyxFcBPChF1w9w
EPD1J/cMaucGhHlxt/DZQLT13RHEMOoSesHbVgntXq3fgGrFdsnmQBtVNxdne99eP8mOErkx+x3+
wgQGE6xPRrYmNVSXqLV3Lr3h9WXYPLedMXS5/xGSRdLeKGAbGMVAFt6X9V5A+a8sjcs3D56sZ4Lz
T5UNoPh0xTAyokylvr6HPYJL3Z22Xrw0fENZBGSqHGPGPmOtY3IfACuY3OdoEPy/49uvS8kJ1sld
NqORY24FHIVX3cbu+MxB8Hybm2RM5sKc9zo9mnpEowYh0Rp/tkyzulyxcF4HC6qMdl2BpqvxSqas
lWBtBStA9ftm/8oqsyyYnKz4tJjwPu7H8vgjZCrePVcLV3KllEbzR6w9OEfiBDqEJOHhrL0VJrw4
2WcRYpajOfwnloDkA3FWKqtjz1xameV4+wi7F2lmoFz02TP1s9HysAxijfwIyaJRlGA14AdmfPZv
q8mDJRD2F3LBA9MpWMBEsf1jYpUEXSO0ec3X9HUhJajOnJE8NYJaRYhh7m2thwTMag6nGkYFfUyO
LpeqiGbq2H0RigMajyHu5OOoPin33lnM0oyntobin3fj+I+YMnP7u+wSaV5R6qgeFSZXdO5aphKk
QidngT9eYXWTRLZoL/75KqzRXjTmqDVVq4YHZRyLOwudg+kISOaT0Wh3/KI5peVPKJ8UdbT84jUn
G4cVVt6Egul3sZIvUewpWBU1MovwtF1UZdijmg//peWCg1msjsd7ztdijhNCh8XoMhMd7RTTesYl
/d2ZSDSzDxt4e+hZNCX3Lqt6ipL2aD0zGXcicBVBnKt0POs/xnLnkuiHSY7+IGoysCufwjdn8qRl
X9eeGwMEPlZcMBvx6wuvV982zxtRamvfFfN9e+4XhRkVYH2AzbgqjCMTngxDYOVlaTq98xgl3B5N
b3S+Si1ndd3K3wCol4hh3GGIWR6IEPKmGSjdK+vfOEViNCu5L4fj/lByHFTZzUiIde+7t6oAyNM4
ii4XEdOzqw4K9wyv80J2D5hHn+YFqdodZbm2I2Sb2ujHdlFeEW1N/0MDeZ/aorhyGbGh3wosRDBa
GYzVs7PiftdXT4d+bS1JpR+RRXMWCF1N6XwTQzzLKjxNmBuk2r1wXsfyLIr6CwpSYVi6Nj1PhAEE
4CaxLJTosQFZig4F4XGlizFfDegroMLyZHhnS2ZtzZNnTnTxG+ir/xU+89iCnozgOt0x1npa/KnJ
jUQAaWik3KdJ8rmt3+4Jm/R3zhRzFFFqYfstd4KVsbbJ5PduPs54i6pjnF+IkOZIojCeqN2a0zIX
ByRGCj/R1LrkKGUtBNQHzIEJ8mQJrvgv7sx2bNjxvA5u4y3jK50rIlwCpVIRGGnE2wIcnoZQaSwD
f8HVgYc+aRqCTNXttu6NjoqaRfgiB2DLjbdcVGyDaGe/5RdhDM/KHtuMCkF7bW9R5Laur+ueBCJK
Q3RwgQNsmDDyE8zy1NxCCZk2BnU4tNUFnfQpFXabUqDykOmrxo9X/WEut/vSJOaAD0tgwY2oE2AO
66MCRE9NqIhaz/ujEh24XaSdb00WfIiqCa9kXhyCMSO+R87kkqT9KkJ1mxTUZItDFHVnD7sFsqCx
O88nm/ycA7MKr33SlB0SXeCii7zILqWVKV0767u9oqI6xvEk/2jmeY2iIfnmkMEx9CKDMwhM3rwu
zoagHMKhRnbF+oich8cpk5uyTPfZt264yyHgs2cbrOOomrUXPw5lBT+66kRwCwWs6GN6XZHQz2Dg
uZwR0DgTHr4tI1wmEWOTiWg/0wRJgD1C2azKPakLNGb4s3WuHWpF5COizMJyqrwtjb0pRarmQ/mD
SLCHNmWVzHGEXcJ2gURHsZnNUK+Ibq99c9rBfoIf56P1KWkTGIbVTeZNHMXle0G0A0wK1DiiENs1
T4IuF67PPrZ9TFs9lpSI/bkyPLdWb15egKMBfNOmnKHqZJ6B5xmDARqG2eE8tZtX41JGMkd/fNf+
Bw+gpoMP9p51SlrpNp0WozW6uiD0qvtKQ0lKbAGmWG/nDwejpItLVb1j78bXcjVHK23gsKzoO3yp
4LuEUXBva8Q7on5H0bVjsW0v5YC3wrv7filttqLtsxGF1PIG2BSYnCIMMv1kzy7Nq5rxZboXXL61
Hkkwkbk3Zoy7ZtA3aPaEUZX8YdCtaIYxlNx51MkaX08I+huCwAHR7XaqdKHZJI+cXRk8goz0H38K
dCRrBcTC4IJsexHsLgnOqFOJ+lIPl2URlsKLUB9rRrnjRwHfjWM16X/f+cVj0ppVoaIyQxqkkOLr
eUh7mJHkl0/Kw2fVzD4E3MzbHhpkGTVVYl8Ep5vP7bcAfIt/Ixmp82wRB14Dr0VwK+4dy/51K27s
IY7vcOHAdeIf/YDj6+XhIxnfyZv17XKZ+NPrNHB6+osJRjCH0fAYfWps7Idax0q2562l7RU0Nmnw
AjFYMoY7KS83jDNqFc8zxwSehindljxlupoKjG4v86MXLInPWB/lgYxczV8W6i0LPL/k777ZDs6K
F0NjMoQ4UYOXc5rho39zKdVXtTuD/vRgcb4R3CmdlpbxOkSbir5IvQURqV+RdwWKrwFILKaI4K5g
Z2tjhq3KSRVDvcJatmVYwFMjbiYW4ydmLpjSfeQZyTkhP8Kpv2F0YAIETLO4uL5CxaO8zvVtxnLY
BsJji4KseMb5mDY3CL3TUUN1bUquimtW6ceUo5ReseBL/R586d+Q2wXWyPb4jycfNHWgOcYR8iWE
8YCL7Z6GjeVcRUMfrBkRdUpthn5WESZTD4pfaF60T8Fhj0sHNpUeGckBwdPRzB1YxTO5H4pWBmoC
ZSO+pBibjMq8+czcbjSzcM8whHkf0O/BOamf2Tg/zgS8BvXQhA8lwFmYhAjugWXQlKL65j/53mSH
wXFpmhtyjAp6HtdfSvhWY/OT/3F1fMBE1HDBFU9d+rkKfNBhcnu2SAKsuTEuSRdnm2jYpPVU09xC
093vDUA+LvHNfEX1KEUk/K6hqcPzZyIdNinAiQjsNeQM8tNc1FBttjXy8U5ZQrbE1aSuCNq8BDKI
LZCEpkbiuixqC+BS6lCo+wC9u+w4yjx2k8wI9E9QDpypDKpUgq84+hljaHUbUuJUEcnPLgNXEAX/
riix8tQr1z9lHC9gr3yuJiWa9/7ewak2yowKEXwRMxJvWvntDJYMcgo1hhfS8GSNBMjcRLQWeg7L
iRnpiRIo9oEuhPUhPU1MTGhJpRiSMeTqErgjDw20bDsUaPqd7B7sZ3rsomSwQu4vi6JD/D3w6xKE
GGo+7QU1ECzKk0/tfhzsCmTcjCaO8MFVafSJXJzaE0f88kofm0k7zeWYcl3Ns1vqnSYISSfBzu7Y
B1HxsB16M3efuaG3UEv1F7l5UgPAA9K42zRx2rIn1LEy6tI4SZDtJprAouKVkPQ6spoRJwiGyzxw
j5xouC1jmmbau4uVlEQH/wKRjUDohEMBxNX1P3IkjcLSMraHx0gnZI0NfDZ/ldA96fOkfafPAjdD
5h3u3xynegUvFeql4K1urhmPLVBZjQq2Q9mwtBfmyDb8Q3rvbd82ulDZ0juVbIHVv2fsL5OzcG5L
IDfm83Dn+dYHeUsUTozAFjKdSP8L6Ci8XDdlCXagvTb+xQXU0m+5y2774Pl7f8TuMoYqNY+8aryT
8hawUwyzNORwX8v9a2O4y1g0aNrqP3sIsBRC366RTsoqrUd7GDxXI93qzRiBkdoC5HwKj2kpI1ee
94JytXIrfIilq3tkJrYpfak/tNKgZlMMtq/N0llJ8QiMDjDhNpLAYnGdScLB0laspFyWSjGmD6ua
yCjIPfSB+mK6Srkp5QbiQElnDpYQO0Q6umNyA5RcEyJswarRMeMaCrzhjqz9KP1Q+2F9QNpltOOr
Llcm82F/7XdQjlIU1WuvyrogDrHn/ffN9dH0dyis1sn2wyPl/bDvgnbqZUDo2h1JOF9Nh9IA/pLk
6MJ0L35iF8toNv+NAUprDE8pIfLAe5vRypf5gnH9VNZkoKatfnJh5ztEbLxOpovex+QGsY6f7oWS
g/7+MzfVGuFEy4+hXK44vjV6vrFPpvDSYEImqFMFitCGouaADyNM+RFjavFH1EVToFqkoYcGxudj
HORzMzG4cduR2mhYS5vUhZHJ81FOowlLr4rpdeIBrVarEsPFLbWsALgnoH0X5bkxEF4E0A268z72
kDkELelh4Nfv5e+TTeIMxTMV/H1knWvs3JO8XTRi1AKlzYqJpMYTkSO1o8mT6jx4JYi4RrfNtR5o
QPobcTl7uIcppoTEwcjmSYUcTIvsQn+Ax0X/5uNCss8Kuz2vYKeRrBijCnpppY4TwWLQJrYkF596
aOZiYuuY5vCNSzWoWp7uve72xSqYwenHdWpvt2/Ggrq8D+lhO3R5WtYfLFoMmoy/CYGgG8Iixio+
Vjcbl1BQy9zLEzchXs+v95YZcATV/bwq/2LKgtfMm5c0O8OhgM/OZJU8efrRiNGf5O/0YUO/Oawg
o2LBloe2C4vHR6Pg8Wu8D1V/CHXfAZVTqrMWiMKDdmE4zAwD2xyCmsPi/Ycf69Ch7kT8ZaCxiBKj
CfHT11YVjwsZ7rGJtnMvlD4UICeoqvwZ/Gw/Tnm48hOmnJrvHf0ryG8b2mG5TyJi3XjyIRS52qw/
grDoUwF/IFZ+PeRCtqDr5PqT5yx/qI3CYCwxL9NoiImrSRCDfx0LaXFyhlyMlC49YOqXilyLTJGp
4wp9//hene3rPLQyxpb9Ug5wDiz36GINj679GOsYV3nWiUr6ibWLqAjAO2AiQZzQyWpznnG1Nz4d
VmBG1j+3sfYPLvWXPtuWldA5zO/yMGJolqVElx2+qnGyi+m3G+6Oj5yoN+V3HEZLbGgHWJQnj1QN
tqvH8KNR13k/kBqdi2w5kUP+TMlfQ9fEd1LEbccW7F+Rw2N91721/nf1Y0gszITVm8Q3r1libKvK
lbIZwquu/hPwtskTdXXhN2YfhI0W6LF+T6KUhc//d6FZCvGpaeWbbfoUVMccm2QgQJS0jUTvs6ad
Zr4SHcTZx1Pd4BFIH+rmYmlJ4emTjTeO4ZB+t5wSk+YmChx9/Aw27XmNcpLJ9xZGJNmDw+wPCPeG
Kf5hLgHOW+liVwis+obFGthQVF/cYfiVNmZM/osSC3YfDBCqjbw8FQOVf+h14dqHqKdbUf4RE1P8
PemvBYvdyqLDg3YMzahO2k0SKKdWd3+MLRf+yZvwcNUSshikSyphJycq4245TRc7yxEuCRs9FH/e
wBmkwYxwvqiwwvVZ5ODNldq4AKgCM5ANo4OCbI+k+Yy5UaZM4rEMYaA6gqMzSEdPouA+v4zgcBjb
CztGgCx6+s8ThVn+CGxfkcMxfFYMUURFrYkUuqCXHRec6IHp8KgNXxg3YvTEP9OXZGTs06KTduAe
xWSbdP0/vwWDN9k4JU/h6NoI1858U1Yu6OnoCFg665Nm9OoaVTuofGh7sM2tt3Ecc8IKPEmdgvqY
v8t4aaxr0JI8IvUBITBwRv2RxGwosxI+x+KSCT2gav2zzL67F4Gw7ftA1JSy5OotsajaBZw4Qqlc
9LTZNwFASmk7UsxykstaLAN7jhpY0zyw/i190OfnUKBOaEnNkiRLEfNYIEU1ZR4i73t/64sSbWkQ
5YxjLtqTKbVMfFv/8jf/VQ7Vj4WT2OQSjYy0xZexKhZWRJAyCHZJHzuXfGvJK0avGYpALDpmveCG
tused4tbMePMaAFHJIwxLjRNu7JngZk7eswLxd8X9EKQeiqblCWbJOS/cGHt4i72cKpN7EsZYrR2
iCStMSxg2JOy0QQymu/1hiuHc+5rZ6KUIVsyCUkFQah/3h7Evvaj3kTonk/yMrVhS2gC9hpsC3Vj
Sw/6C1lBIjJOGiTd0VAXcvkuElbu0re8nUEHENAd3CaeEbtcmr0Hn7WUFaIWPZ0jvrlSJLUPVf/D
f/2kkciAoxNJvSS5VDfEeg22q6y5/woJijV6LpqYUhLBk+Hggcd4pWPNpAd3HBlLuRtVX7SeSgTr
Aj5NaHtuhueBKFihlyhjkMKmAEKG3hMTAicHCJt927DW+gC6Uhiibq/6yW4rAS2dtyxbc8wjtZIG
VO0XDL0QdvxkJ4/ihMj36blL/07MQiI8SmrW16ItX8zBYfgyiPnKTVTlbWmbnGwQz0RuQjUmuDi6
xWBriT3wIcoi6iriQ09fqcK9yJEKsjZRfa01Bf8XG+iP2EqZjE/BaAqLoHeQE6PGhn5Jlaxamx5K
rMG426GbTw8QHam25GhDobv9sShlNmr0EJ8kFZL3tFZYC7HtZNyzG572L4alFxA5pf9gPOeuq0cg
Kfss0Tn66Pr7ONw/Iu6uVVaMsfkRFy4gVPZhv40c8nd0P0nlVUbM4NiYvHfKKh+1ULstT3RVr6U6
7994y373xcsMLvC/M8F7rJprHNIHFLb2EG5WBTgK/p8xzDvzF09IriuqH+QmqoKCYdpDmWLLbOV+
WbhMMvb230vxUeOkgz0J8SJfRx5SBJ1TfoRVPyeGhX0VCH0WWSLRXJNpSC6cPijEwx0YBkF96s69
Yn7ILlCVQJxLD6WmDzfD1193GYLWLtoeB7OXVThM/bxgIG3v2H0z0TAOOPI/c2awY1RPJTuhMiB/
HOl9RS9iustYPGt29a8MOk3hqkzKct8xQQG1nl6cnU5PWOQGA+yCco/HMvSKBGOqXYBsRZ5N2Auu
7ZME3nmGmHOXm/h0hP85kuUKENpTpn9+cSQTr1feRH+BbCtc1l1g65T/ahtx0aEBmIdrk3a/wZJq
JHVPiczz9B/B61Kn44jcB3q/DJxcnzoyZAvWq6bwuWEy06aCwNL7zcVR28LTfE2Lxwj4E0jcY1Bh
aFX1pmuPw9D3xC2YCwLAf1Td8VYfafXdL+08oNiiRsnnI6ZtetKlu6jMnEHi30EVC3OOvRGirjv2
tbzkr3bgGTdJddvGF5+hOkJavUs1c/YfscBgdZvA5gZ5fPfknkPjlV0KzvBHngyq6wig9zE1QwJN
e9M+08NpcBxN5GdDtImaoJhSi8EqS9nxqi4P3zanFcrZ3l0JuZJ2QHACRDT4JioleRJ0maSHC4cz
mRALZjtwWfI+iH4qtR/Hqz3rgF55hlCj1yQNN9NfemWFnJBu0UVuw1uWgG0+bHu4vcHfZpRwP06W
0pr/a1bFXIdQI/AXa1hBruYuXNnVL+jAm7MlnPkp8Zn0qU74NCAzGUkxFd24RRQjcWzkcj36h1HJ
JOTXU/igTvr5hzd/w0ms3bvj+V2PI7Heb1TxYGXWuQMicP+G2e7KtsMKjX+BH7qeNt0I8Spc4jIM
ATX7QttN9geQVceI0SW7QTbHnAX7fJKC2M8fwOV6GEGrr4X5n4oKDi7qGxg5uhtmBu1XPtF+pApp
vpoxtR4NnUOo/VnEFGumxyYJhK6r+TEx5OA78aDmXV+tuhdC6pMMaI+9e66g0iqvoGOPOWlfly+h
0cXFxyQO7kHmJQ8sSK/4OOpGeOaDyDjejj8jSaKu4ducEgGuOo9gWT8GmW8G+oCcwoCIcBn7iNfJ
oLJyukharrhfW1apNupzaTOjoOPknsCDaVUm6jCEBpJzF1Nm9208id10XRh3TJpj45Jw3T+HPwel
38gVNdT1znD+PTD1ZCa66BMw3pDCkBybf+sZRQppmtee2jcn2cKyPk2gHus7covza0njMXWi8X4+
+ZmIgzA9j6X6o4clfiWGrUwOYWvtw5lQVUNTShrEnO5LKhFhP6Lp+o3Np1skqwRjQKP1ls1gCXJq
MaDw6sbMb5fX/QFObVbSzKU/tgocEXfVBgJSNgNJGg1lfI4y9VhvwbssdCxKMtJPvtxnH7/r7nbX
Iw3qJu5kmRfHcec7gqo7XGW7JGzO44l2Qv7lLCu1sf385yvhu5CT3vp0JztswHnHHxZes1htZs5A
TUYpnrgIxJUjd5BQoZb7m3Pt9PuKabOWdlw7QalX3FTwe/Sc0gVL49er70KDM7tlgOUFNkSSXzM5
oYI9mc3I4kfUWL/gO/nfebcEmAOEheO8NGRSZfdtXzNj9sRoCnd7+zCobhFFh3rkEJIiGTksXpcI
CQOnB9fCsiB21RYc6/8yAPHUP2lU4an2WNZbYxd5rC9R4dVnvoPZJmZFi9aX9X3goVnaC3FYPddk
g5b/JITnbQmPXDXbVb3Hcg7Ep8iPkhthAzNeudN8sHcp6Oc81D1rhgtcRAM3fC2pjMVLYLNDs0fb
MGl1y+CLIz22HnRIbDEX1tlJvvqnVmRpIffHPKh4zjzHO+VOrn/gdjTrSQ1cAuwTy48OlVFMKZ3n
fgnMk+I0Q77+DwebCHsoTTnKjRGnk4Jq6uPsWOrHr5RsJ75AjI9YrtUtC94bq5Y2UQm9OhizhiSG
iNda/dTHS31j2s/4aSgEdT6nxm+ptsPs7haefxvJroT8f9uHLIgyvKPcEKsYL7knssNwtz4nHxjo
cfG5hg67zy1NM/3BqbmEvgUd8bs1kFBUEEFcxZvlL24y4mSSPoTX21y7Nv3e1rafSuHFCx8l6zIO
1hIseYWChWSFoGXr/AS98fXBFI7HBHGT1biBMZ5Tb0ot2x8jScIj8sHlinSOTsT6mWBpTj4uHTEg
Yd9AWbrqjw7yuYNCzT7tfYFMKbD65EePm45DhPyYDeKYSCALwuXCTMfXTRyHN0GHf7/TWmlSUOPG
YsTid3AuFd4+X2dOo8u8pQ2w20e2VxEJWbR7csZY7KKaUah5AfOIj3XDuyMr83azjx/76325nTue
XswKYhHPYmSrgksLKiNOHpCLAMH/luJMjStUxfd5g2V6kykxqxM1fs0DR9u9Mvw83bYMR6qgjse/
/0Zcqu6bqjOF6q5HjtG5G4o7m6z/foe72i0eaAU2GOmZLIO1SDOIcPgSxr5cuZUW5ieevziGv6UI
g+kNLR4F0fOADyaX/gPKBbxwgaO/BwQehGNqhxftK11ce4BAQFYGH+hpOGyHC2tUzERaLqcQsBRS
sM48GZ5VVVFntw+2+upaGKb2VaFYTW11c8xhPe9DSarWsk3MeKhfS7be0AplOXcLjFC4G3ldsiXv
AgAETvoJstGfVrbucsT3QpTLKPcf75HPBvamokDSUklv4vG3UJwJj/+MBYtmN9pXYAmPiHfWUjjT
DvKnat+wowx/KD+ukpQ5UGglTuh/Nsoueeixdc3aHO/YtpJ0093W4/X1itcOzi1HoVwmGnAGn8R7
SpLelqYURdXyp2Z1rdaNyTqztv7vaLTNu6/hOMO26R2rIwometHW51EgLJ0IsIzsu6+KQo2KvbSX
1OO9dzyPZEA8eFu87hAn7gvlJFB0bw==
`protect end_protected
